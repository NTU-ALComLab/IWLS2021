module Conv22(
input [4:0] x0 ,
input [4:0] x1 ,
input [4:0] x2 ,
input [4:0] x3 ,
input [4:0] x4 ,
input [4:0] x5 ,
input [4:0] x6 ,
input [4:0] x7 ,
input [4:0] x8 ,
input [4:0] x9 ,
input [4:0] x10 ,
input [4:0] x11 ,
input [4:0] x12 ,
input [4:0] x13 ,
input [4:0] x14 ,
input [4:0] x15 ,
input [4:0] x16 ,
input [4:0] x17 ,
input [4:0] x18 ,
input [4:0] x19 ,
input [4:0] x20 ,
input [4:0] x21 ,
input [4:0] x22 ,
input [4:0] x23 ,
input [4:0] x24 ,
input [4:0] x25 ,
input [4:0] x26 ,
input [4:0] x27 ,
input [4:0] x28 ,
input [4:0] x29 ,
input [4:0] x30 ,
input [4:0] x31 ,
input [4:0] x32 ,
input [4:0] x33 ,
input [4:0] x34 ,
input [4:0] x35 ,
input [4:0] x36 ,
input [4:0] x37 ,
input [4:0] x38 ,
input [4:0] x39 ,
input [4:0] x40 ,
input [4:0] x41 ,
input [4:0] x42 ,
input [4:0] x43 ,
input [4:0] x44 ,
input [4:0] x45 ,
input [4:0] x46 ,
input [4:0] x47 ,
input [4:0] x48 ,
input [4:0] x49 ,
input [4:0] x50 ,
input [4:0] x51 ,
input [4:0] x52 ,
input [4:0] x53 ,
input [4:0] x54 ,
input [4:0] x55 ,
input [4:0] x56 ,
input [4:0] x57 ,
input [4:0] x58 ,
input [4:0] x59 ,
input [4:0] x60 ,
input [4:0] x61 ,
input [4:0] x62 ,
input [4:0] x63 ,
input [4:0] x64 ,
input [4:0] x65 ,
input [4:0] x66 ,
input [4:0] x67 ,
input [4:0] x68 ,
input [4:0] x69 ,
input [4:0] x70 ,
input [4:0] x71 ,
input [4:0] x72 ,
input [4:0] x73 ,
input [4:0] x74 ,
input [4:0] x75 ,
input [4:0] x76 ,
input [4:0] x77 ,
input [4:0] x78 ,
input [4:0] x79 ,
input [4:0] x80 ,
input [4:0] x81 ,
input [4:0] x82 ,
input [4:0] x83 ,
input [4:0] x84 ,
input [4:0] x85 ,
input [4:0] x86 ,
input [4:0] x87 ,
input [4:0] x88 ,
input [4:0] x89 ,
input [4:0] x90 ,
input [4:0] x91 ,
input [4:0] x92 ,
input [4:0] x93 ,
input [4:0] x94 ,
input [4:0] x95 ,
input [4:0] x96 ,
input [4:0] x97 ,
input [4:0] x98 ,
input [4:0] x99 ,
input [4:0] x100 ,
input [4:0] x101 ,
input [4:0] x102 ,
input [4:0] x103 ,
input [4:0] x104 ,
input [4:0] x105 ,
input [4:0] x106 ,
input [4:0] x107 ,
input [4:0] x108 ,
input [4:0] x109 ,
input [4:0] x110 ,
input [4:0] x111 ,
input [4:0] x112 ,
input [4:0] x113 ,
input [4:0] x114 ,
input [4:0] x115 ,
input [4:0] x116 ,
input [4:0] x117 ,
input [4:0] x118 ,
input [4:0] x119 ,
input [4:0] x120 ,
input [4:0] x121 ,
input [4:0] x122 ,
input [4:0] x123 ,
input [4:0] x124 ,
input [4:0] x125 ,
input [4:0] x126 ,
input [4:0] x127 ,
input [4:0] x128 ,
input [4:0] x129 ,
input [4:0] x130 ,
input [4:0] x131 ,
input [4:0] x132 ,
input [4:0] x133 ,
input [4:0] x134 ,
input [4:0] x135 ,
input [4:0] x136 ,
input [4:0] x137 ,
input [4:0] x138 ,
input [4:0] x139 ,
input [4:0] x140 ,
input [4:0] x141 ,
input [4:0] x142 ,
input [4:0] x143 ,
input [4:0] x144 ,
input [4:0] x145 ,
input [4:0] x146 ,
input [4:0] x147 ,
input [4:0] x148 ,
input [4:0] x149 ,
input [4:0] x150 ,
input [4:0] x151 ,
input [4:0] x152 ,
input [4:0] x153 ,
input [4:0] x154 ,
input [4:0] x155 ,
input [4:0] x156 ,
input [4:0] x157 ,
input [4:0] x158 ,
input [4:0] x159 ,
input [4:0] x160 ,
input [4:0] x161 ,
input [4:0] x162 ,
input [4:0] x163 ,
input [4:0] x164 ,
input [4:0] x165 ,
input [4:0] x166 ,
input [4:0] x167 ,
input [4:0] x168 ,
input [4:0] x169 ,
input [4:0] x170 ,
input [4:0] x171 ,
input [4:0] x172 ,
input [4:0] x173 ,
input [4:0] x174 ,
input [4:0] x175 ,
input [4:0] x176 ,
input [4:0] x177 ,
input [4:0] x178 ,
input [4:0] x179 ,
input [4:0] x180 ,
input [4:0] x181 ,
input [4:0] x182 ,
input [4:0] x183 ,
input [4:0] x184 ,
input [4:0] x185 ,
input [4:0] x186 ,
input [4:0] x187 ,
input [4:0] x188 ,
input [4:0] x189 ,
input [4:0] x190 ,
input [4:0] x191 ,
input [4:0] x192 ,
input [4:0] x193 ,
input [4:0] x194 ,
input [4:0] x195 ,
input [4:0] x196 ,
input [4:0] x197 ,
input [4:0] x198 ,
input [4:0] x199 ,
input [4:0] x200 ,
input [4:0] x201 ,
input [4:0] x202 ,
input [4:0] x203 ,
input [4:0] x204 ,
input [4:0] x205 ,
input [4:0] x206 ,
input [4:0] x207 ,
input [4:0] x208 ,
input [4:0] x209 ,
input [4:0] x210 ,
input [4:0] x211 ,
input [4:0] x212 ,
input [4:0] x213 ,
input [4:0] x214 ,
input [4:0] x215 ,
input [4:0] x216 ,
input [4:0] x217 ,
input [4:0] x218 ,
input [4:0] x219 ,
input [4:0] x220 ,
input [4:0] x221 ,
input [4:0] x222 ,
input [4:0] x223 ,
input [4:0] x224 ,
input [4:0] x225 ,
input [4:0] x226 ,
input [4:0] x227 ,
input [4:0] x228 ,
input [4:0] x229 ,
input [4:0] x230 ,
input [4:0] x231 ,
input [4:0] x232 ,
input [4:0] x233 ,
input [4:0] x234 ,
input [4:0] x235 ,
input [4:0] x236 ,
input [4:0] x237 ,
input [4:0] x238 ,
input [4:0] x239 ,
input [4:0] x240 ,
input [4:0] x241 ,
input [4:0] x242 ,
input [4:0] x243 ,
input [4:0] x244 ,
input [4:0] x245 ,
input [4:0] x246 ,
input [4:0] x247 ,
input [4:0] x248 ,
input [4:0] x249 ,
input [4:0] x250 ,
input [4:0] x251 ,
input [4:0] x252 ,
input [4:0] x253 ,
input [4:0] x254 ,
input [4:0] x255 ,
input [4:0] x256 ,
input [4:0] x257 ,
input [4:0] x258 ,
input [4:0] x259 ,
input [4:0] x260 ,
input [4:0] x261 ,
input [4:0] x262 ,
input [4:0] x263 ,
input [4:0] x264 ,
input [4:0] x265 ,
input [4:0] x266 ,
input [4:0] x267 ,
input [4:0] x268 ,
input [4:0] x269 ,
input [4:0] x270 ,
input [4:0] x271 ,
input [4:0] x272 ,
input [4:0] x273 ,
input [4:0] x274 ,
input [4:0] x275 ,
input [4:0] x276 ,
input [4:0] x277 ,
input [4:0] x278 ,
input [4:0] x279 ,
input [4:0] x280 ,
input [4:0] x281 ,
input [4:0] x282 ,
input [4:0] x283 ,
input [4:0] x284 ,
input [4:0] x285 ,
input [4:0] x286 ,
input [4:0] x287 ,
input [4:0] x288 ,
input [4:0] x289 ,
input [4:0] x290 ,
input [4:0] x291 ,
input [4:0] x292 ,
input [4:0] x293 ,
input [4:0] x294 ,
input [4:0] x295 ,
input [4:0] x296 ,
input [4:0] x297 ,
input [4:0] x298 ,
input [4:0] x299 ,
input [4:0] x300 ,
input [4:0] x301 ,
input [4:0] x302 ,
input [4:0] x303 ,
input [4:0] x304 ,
input [4:0] x305 ,
input [4:0] x306 ,
input [4:0] x307 ,
input [4:0] x308 ,
input [4:0] x309 ,
input [4:0] x310 ,
input [4:0] x311 ,
input [4:0] x312 ,
input [4:0] x313 ,
input [4:0] x314 ,
input [4:0] x315 ,
input [4:0] x316 ,
input [4:0] x317 ,
input [4:0] x318 ,
input [4:0] x319 ,
input [4:0] x320 ,
input [4:0] x321 ,
input [4:0] x322 ,
input [4:0] x323 ,
input [4:0] x324 ,
input [4:0] x325 ,
input [4:0] x326 ,
input [4:0] x327 ,
input [4:0] x328 ,
input [4:0] x329 ,
input [4:0] x330 ,
input [4:0] x331 ,
input [4:0] x332 ,
input [4:0] x333 ,
input [4:0] x334 ,
input [4:0] x335 ,
input [4:0] x336 ,
input [4:0] x337 ,
input [4:0] x338 ,
input [4:0] x339 ,
input [4:0] x340 ,
input [4:0] x341 ,
input [4:0] x342 ,
input [4:0] x343 ,
input [4:0] x344 ,
input [4:0] x345 ,
input [4:0] x346 ,
input [4:0] x347 ,
input [4:0] x348 ,
input [4:0] x349 ,
input [4:0] x350 ,
input [4:0] x351 ,
input [4:0] x352 ,
input [4:0] x353 ,
input [4:0] x354 ,
input [4:0] x355 ,
input [4:0] x356 ,
input [4:0] x357 ,
input [4:0] x358 ,
input [4:0] x359 ,
input [4:0] x360 ,
input [4:0] x361 ,
input [4:0] x362 ,
input [4:0] x363 ,
input [4:0] x364 ,
input [4:0] x365 ,
input [4:0] x366 ,
input [4:0] x367 ,
input [4:0] x368 ,
input [4:0] x369 ,
input [4:0] x370 ,
input [4:0] x371 ,
input [4:0] x372 ,
input [4:0] x373 ,
input [4:0] x374 ,
input [4:0] x375 ,
input [4:0] x376 ,
input [4:0] x377 ,
input [4:0] x378 ,
input [4:0] x379 ,
input [4:0] x380 ,
input [4:0] x381 ,
input [4:0] x382 ,
input [4:0] x383 ,
output [4:0] y0 ,
output [4:0] y1 ,
output [4:0] y2 ,
output [4:0] y3 ,
output [4:0] y4 ,
output [4:0] y5 ,
output [4:0] y6 ,
output [4:0] y7 ,
output [4:0] y8 ,
output [4:0] y9 ,
output [4:0] y10 ,
output [4:0] y11 ,
output [4:0] y12 ,
output [4:0] y13 ,
output [4:0] y14 ,
output [4:0] y15 ,
output [4:0] y16 ,
output [4:0] y17 ,
output [4:0] y18 ,
output [4:0] y19 ,
output [4:0] y20 ,
output [4:0] y21 ,
output [4:0] y22 ,
output [4:0] y23 ,
output [4:0] y24 ,
output [4:0] y25 ,
output [4:0] y26 ,
output [4:0] y27 ,
output [4:0] y28 ,
output [4:0] y29 ,
output [4:0] y30 ,
output [4:0] y31 ,
output [4:0] y32 ,
output [4:0] y33 ,
output [4:0] y34 ,
output [4:0] y35 ,
output [4:0] y36 ,
output [4:0] y37 ,
output [4:0] y38 ,
output [4:0] y39 ,
output [4:0] y40 ,
output [4:0] y41 ,
output [4:0] y42 ,
output [4:0] y43 ,
output [4:0] y44 ,
output [4:0] y45 ,
output [4:0] y46 ,
output [4:0] y47 ,
output [4:0] y48 ,
output [4:0] y49 ,
output [4:0] y50 ,
output [4:0] y51 ,
output [4:0] y52 ,
output [4:0] y53 ,
output [4:0] y54 ,
output [4:0] y55 ,
output [4:0] y56 ,
output [4:0] y57 ,
output [4:0] y58 ,
output [4:0] y59 ,
output [4:0] y60 ,
output [4:0] y61 ,
output [4:0] y62 ,
output [4:0] y63 ,
output [4:0] y64 ,
output [4:0] y65 ,
output [4:0] y66 ,
output [4:0] y67 ,
output [4:0] y68 ,
output [4:0] y69 ,
output [4:0] y70 ,
output [4:0] y71 ,
output [4:0] y72 ,
output [4:0] y73 ,
output [4:0] y74 ,
output [4:0] y75 ,
output [4:0] y76 ,
output [4:0] y77 ,
output [4:0] y78 ,
output [4:0] y79 ,
output [4:0] y80 ,
output [4:0] y81 ,
output [4:0] y82 ,
output [4:0] y83 ,
output [4:0] y84 ,
output [4:0] y85 ,
output [4:0] y86 ,
output [4:0] y87 ,
output [4:0] y88 ,
output [4:0] y89 ,
output [4:0] y90 ,
output [4:0] y91 ,
output [4:0] y92 ,
output [4:0] y93 ,
output [4:0] y94 ,
output [4:0] y95 ,
output [4:0] y96 ,
output [4:0] y97 ,
output [4:0] y98 ,
output [4:0] y99 ,
output [4:0] y100 ,
output [4:0] y101 ,
output [4:0] y102 ,
output [4:0] y103 ,
output [4:0] y104 ,
output [4:0] y105 ,
output [4:0] y106 ,
output [4:0] y107 ,
output [4:0] y108 ,
output [4:0] y109 ,
output [4:0] y110 ,
output [4:0] y111 ,
output [4:0] y112 ,
output [4:0] y113 ,
output [4:0] y114 ,
output [4:0] y115 ,
output [4:0] y116 ,
output [4:0] y117 ,
output [4:0] y118 ,
output [4:0] y119 ,
output [4:0] y120 ,
output [4:0] y121 ,
output [4:0] y122 ,
output [4:0] y123 ,
output [4:0] y124 ,
output [4:0] y125 ,
output [4:0] y126 ,
output [4:0] y127 ,
output [4:0] y128 ,
output [4:0] y129 ,
output [4:0] y130 ,
output [4:0] y131 ,
output [4:0] y132 ,
output [4:0] y133 ,
output [4:0] y134 ,
output [4:0] y135 ,
output [4:0] y136 ,
output [4:0] y137 ,
output [4:0] y138 ,
output [4:0] y139 ,
output [4:0] y140 ,
output [4:0] y141 ,
output [4:0] y142 ,
output [4:0] y143 ,
output [4:0] y144 ,
output [4:0] y145 ,
output [4:0] y146 ,
output [4:0] y147 ,
output [4:0] y148 ,
output [4:0] y149 ,
output [4:0] y150 ,
output [4:0] y151 ,
output [4:0] y152 ,
output [4:0] y153 ,
output [4:0] y154 ,
output [4:0] y155 ,
output [4:0] y156 ,
output [4:0] y157 ,
output [4:0] y158 ,
output [4:0] y159 ,
output [4:0] y160 ,
output [4:0] y161 ,
output [4:0] y162 ,
output [4:0] y163 ,
output [4:0] y164 ,
output [4:0] y165 ,
output [4:0] y166 ,
output [4:0] y167 ,
output [4:0] y168 ,
output [4:0] y169 ,
output [4:0] y170 ,
output [4:0] y171 ,
output [4:0] y172 ,
output [4:0] y173 ,
output [4:0] y174 ,
output [4:0] y175 ,
output [4:0] y176 ,
output [4:0] y177 ,
output [4:0] y178 ,
output [4:0] y179 ,
output [4:0] y180 ,
output [4:0] y181 ,
output [4:0] y182 ,
output [4:0] y183 ,
output [4:0] y184 ,
output [4:0] y185 ,
output [4:0] y186 ,
output [4:0] y187 ,
output [4:0] y188 ,
output [4:0] y189 ,
output [4:0] y190 ,
output [4:0] y191 ,
output [4:0] y192 ,
output [4:0] y193 ,
output [4:0] y194 ,
output [4:0] y195 ,
output [4:0] y196 ,
output [4:0] y197 ,
output [4:0] y198 ,
output [4:0] y199 ,
output [4:0] y200 ,
output [4:0] y201 ,
output [4:0] y202 ,
output [4:0] y203 ,
output [4:0] y204 ,
output [4:0] y205 ,
output [4:0] y206 ,
output [4:0] y207 
);
wire [13:0] sharing0;
wire [13:0] sharing1;
wire [13:0] sharing2;
wire [13:0] sharing3;
wire [13:0] sharing4;
wire [13:0] sharing5;
wire [13:0] sharing6;
wire [13:0] sharing7;
wire [13:0] sharing8;
wire [13:0] sharing9;
wire [13:0] sharing10;
wire [13:0] sharing11;
wire [13:0] sharing12;
wire [13:0] sharing13;
wire [13:0] sharing14;
wire [13:0] sharing15;
wire [13:0] sharing16;
wire [13:0] sharing17;
wire [13:0] sharing18;
wire [13:0] sharing19;
wire [13:0] sharing20;
wire [13:0] sharing21;
wire [13:0] sharing22;
wire [13:0] sharing23;
wire [13:0] sharing24;
wire [13:0] sharing25;
wire [13:0] sharing26;
wire [13:0] sharing27;
wire [13:0] sharing28;
wire [13:0] sharing29;
wire [13:0] sharing30;
wire [13:0] sharing31;
wire [13:0] sharing32;
wire [13:0] sharing33;
wire [13:0] sharing34;
wire [13:0] sharing35;
wire [13:0] sharing36;
wire [13:0] sharing37;
wire [13:0] sharing38;
wire [13:0] sharing39;
wire [13:0] sharing40;
wire [13:0] sharing41;
wire [13:0] sharing42;
wire [13:0] sharing43;
wire [13:0] sharing44;
wire [13:0] sharing45;
wire [13:0] sharing46;
wire [13:0] sharing47;
wire [13:0] sharing48;
wire [13:0] sharing49;
wire [13:0] sharing50;
wire [13:0] sharing51;
wire [13:0] sharing52;
wire [13:0] sharing53;
wire [13:0] sharing54;
wire [13:0] sharing55;
wire [13:0] sharing56;
wire [13:0] sharing57;
wire [13:0] sharing58;
wire [13:0] sharing59;
wire [13:0] sharing60;
wire [13:0] sharing61;
wire [13:0] sharing62;
wire [13:0] sharing63;
wire [13:0] sharing64;
wire [13:0] sharing65;
wire [13:0] sharing66;
wire [13:0] sharing67;
wire [13:0] sharing68;
wire [13:0] sharing69;
wire [13:0] sharing70;
wire [13:0] sharing71;
wire [13:0] sharing72;
wire [13:0] sharing73;
wire [13:0] sharing74;
wire [13:0] sharing75;
wire [13:0] sharing76;
wire [13:0] sharing77;
wire [13:0] sharing78;
wire [13:0] sharing79;
wire [13:0] sharing80;
wire [13:0] sharing81;
wire [13:0] sharing82;
wire [13:0] sharing83;
wire [13:0] sharing84;
wire [13:0] sharing85;
wire [13:0] sharing86;
wire [13:0] sharing87;
wire [13:0] sharing88;
wire [13:0] sharing89;
wire [13:0] sharing90;
wire [13:0] sharing91;
wire [13:0] sharing92;
wire [13:0] sharing93;
wire [13:0] sharing94;
wire [13:0] sharing95;
wire [13:0] sharing96;
wire [13:0] sharing97;
wire [13:0] sharing98;
wire [13:0] sharing99;
wire [13:0] sharing100;
wire [13:0] sharing101;
wire [13:0] sharing102;
wire [13:0] sharing103;
wire [13:0] sharing104;
wire [13:0] sharing105;
wire [13:0] sharing106;
wire [13:0] sharing107;
wire [13:0] sharing108;
wire [13:0] sharing109;
wire [13:0] sharing110;
wire [13:0] sharing111;
wire [13:0] sharing112;
assign sharing0 = $signed(-{2'b0,x222}<<<3'd1)+$signed({2'b0,x23}<<<3'd1)+$signed({1'b0,x287});
assign sharing1 = $signed(-{2'b0,x248}<<<3'd1)+$signed({2'b0,x49}<<<3'd1)+$signed({1'b0,x313});
assign sharing2 = $signed(-{2'b0,x200}<<<3'd1)+$signed({2'b0,x1}<<<3'd1)+$signed({1'b0,x265});
assign sharing3 = $signed({2'b0,x176}<<<3'd1)+$signed({2'b0,x304}<<<3'd1)+$signed({1'b0,x249});
assign sharing4 = $signed(-{1'b0,x233})+$signed(-{2'b0,x160}<<<3'd1)+$signed(-{2'b0,x288}<<<3'd1);
assign sharing5 = $signed(-{2'b0,x218}<<<3'd1)+$signed({2'b0,x19}<<<3'd1)+$signed({1'b0,x283});
assign sharing6 = $signed({2'b0,x206}<<<3'd1)+$signed(-{2'b0,x7}<<<3'd1)+$signed(-{1'b0,x271});
assign sharing7 = $signed(-{2'b0,x178}<<<3'd1)+$signed(-{2'b0,x306}<<<3'd1)+$signed(-{1'b0,x251});
assign sharing8 = $signed(-{2'b0,x254}<<<3'd1)+$signed({2'b0,x55}<<<3'd1)+$signed({1'b0,x319});
assign sharing9 = $signed(-{1'b0,x239})+$signed(-{2'b0,x166}<<<3'd1)+$signed(-{2'b0,x294}<<<3'd1);
assign sharing10 = $signed(-{2'b0,x250}<<<3'd1)+$signed({2'b0,x51}<<<3'd1)+$signed({1'b0,x315});
assign sharing11 = $signed({2'b0,x150}<<<3'd1)+$signed({2'b0,x278}<<<3'd1)+$signed({1'b0,x223});
assign sharing12 = $signed({2'b0,x130}<<<3'd1)+$signed({2'b0,x258}<<<3'd1)+$signed({1'b0,x203});
assign sharing13 = $signed(-{2'b0,x236}<<<3'd1)+$signed({2'b0,x37}<<<3'd1)+$signed({1'b0,x301});
assign sharing14 = $signed(-{2'b0,x148}<<<3'd1)+$signed(-{2'b0,x276}<<<3'd1)+$signed(-{1'b0,x221});
assign sharing15 = $signed(-{2'b0,x232}<<<3'd1)+$signed({2'b0,x33}<<<3'd1)+$signed({1'b0,x297});
assign sharing16 = $signed(-{2'b0,x202}<<<3'd1)+$signed({2'b0,x3}<<<3'd1)+$signed({1'b0,x267});
assign sharing17 = $signed(-{2'b0,x220}<<<3'd1)+$signed({2'b0,x21}<<<3'd1)+$signed({1'b0,x285});
assign sharing18 = $signed({2'b0,x238}<<<3'd1)+$signed(-{2'b0,x39}<<<3'd1)+$signed(-{1'b0,x303});
assign sharing19 = $signed(-{2'b0,x132}<<<3'd1)+$signed(-{2'b0,x260}<<<3'd1)+$signed(-{1'b0,x205});
assign sharing20 = $signed(-{2'b0,x216}<<<3'd1)+$signed({2'b0,x17}<<<3'd1)+$signed({1'b0,x281});
assign sharing21 = $signed(-{1'b0,x201});
assign sharing22 = $signed(-{3'b0,x328}<<<3'd2)+$signed({2'b0,x200}<<<3'd1)+$signed({1'b0,x192})+$signed(-{1'b0,x137});
assign sharing23 = $signed({2'b0,x182}<<<3'd1)+$signed({2'b0,x310}<<<3'd1)+$signed({1'b0,x255});
assign sharing24 = $signed(-{2'b0,x146}<<<3'd1)+$signed(-{2'b0,x274}<<<3'd1)+$signed(-{1'b0,x219});
assign sharing25 = $signed(-{2'b0,x134}<<<3'd1)+$signed(-{2'b0,x262}<<<3'd1)+$signed(-{1'b0,x207});
assign sharing26 = $signed(-{2'b0,x180}<<<3'd1)+$signed(-{2'b0,x308}<<<3'd1)+$signed(-{1'b0,x253});
assign sharing27 = $signed({2'b0,x144}<<<3'd1)+$signed({2'b0,x272}<<<3'd1)+$signed({1'b0,x217});
assign sharing28 = $signed({1'b0,x235})+$signed({2'b0,x162}<<<3'd1)+$signed({2'b0,x290}<<<3'd1);
assign sharing29 = $signed(-{2'b0,x234}<<<3'd1)+$signed({2'b0,x35}<<<3'd1)+$signed({1'b0,x299});
assign sharing30 = $signed(-{2'b0,x252}<<<3'd1)+$signed({2'b0,x53}<<<3'd1)+$signed({1'b0,x317});
assign sharing31 = $signed(-{2'b0,x204}<<<3'd1)+$signed({2'b0,x5}<<<3'd1)+$signed({1'b0,x269});
assign sharing32 = $signed(-{1'b0,x237})+$signed(-{2'b0,x164}<<<3'd1)+$signed(-{2'b0,x292}<<<3'd1);
assign sharing33 = $signed(-{1'b0,x231})+$signed({2'b0,x294}<<<3'd1)+$signed(-{3'b0,x359}<<<3'd2)+$signed(-{1'b0,x103});
assign sharing34 = $signed({2'b0,x310}<<<3'd1)+$signed(-{1'b0,x247})+$signed(-{3'b0,x375}<<<3'd2)+$signed(-{1'b0,x119});
assign sharing35 = $signed(-{1'b0,x225})+$signed({2'b0,x288}<<<3'd1)+$signed(-{3'b0,x353}<<<3'd2)+$signed(-{1'b0,x97});
assign sharing36 = $signed({2'b0,x306}<<<3'd1)+$signed(-{1'b0,x243})+$signed(-{3'b0,x371}<<<3'd2)+$signed(-{1'b0,x115});
assign sharing37 = $signed({2'b0,x258}<<<3'd1)+$signed(-{1'b0,x195})+$signed(-{3'b0,x323}<<<3'd2)+$signed(-{1'b0,x67});
assign sharing38 = $signed({2'b0,x276}<<<3'd1)+$signed(-{3'b0,x341}<<<3'd2)+$signed(-{1'b0,x213})+$signed(-{1'b0,x85});
assign sharing39 = $signed({2'b0,x272}<<<3'd1)+$signed(-{3'b0,x337}<<<3'd2)+$signed(-{1'b0,x209})+$signed(-{1'b0,x81});
assign sharing40 = $signed({2'b0,x260}<<<3'd1)+$signed(-{1'b0,x197})+$signed(-{3'b0,x325}<<<3'd2)+$signed(-{1'b0,x69});
assign sharing41 = $signed({2'b0,x308}<<<3'd1)+$signed(-{1'b0,x245})+$signed(-{3'b0,x373}<<<3'd2)+$signed(-{1'b0,x117});
assign sharing42 = $signed({2'b0,x304}<<<3'd1)+$signed(-{1'b0,x241})+$signed(-{3'b0,x369}<<<3'd2)+$signed(-{1'b0,x113});
assign sharing43 = $signed(-{1'b0,x227})+$signed({2'b0,x290}<<<3'd1)+$signed(-{3'b0,x355}<<<3'd2)+$signed(-{1'b0,x99});
assign sharing44 = $signed({2'b0,x278}<<<3'd1)+$signed(-{3'b0,x343}<<<3'd2)+$signed(-{1'b0,x215})+$signed(-{1'b0,x87});
assign sharing45 = $signed({2'b0,x256}<<<3'd1)+$signed(-{1'b0,x193})+$signed(-{3'b0,x321}<<<3'd2)+$signed(-{1'b0,x65});
assign sharing46 = $signed({2'b0,x274}<<<3'd1)+$signed(-{3'b0,x339}<<<3'd2)+$signed(-{1'b0,x211})+$signed(-{1'b0,x83});
assign sharing47 = $signed(-{1'b0,x229})+$signed({2'b0,x292}<<<3'd1)+$signed(-{3'b0,x357}<<<3'd2)+$signed(-{1'b0,x101});
assign sharing48 = $signed({2'b0,x262}<<<3'd1)+$signed(-{1'b0,x199})+$signed(-{3'b0,x327}<<<3'd2)+$signed(-{1'b0,x71});
assign sharing49 = $signed(-{1'b0,x241})+$signed({1'b0,x240})+$signed(-{1'b0,x120})+$signed(-{1'b0,x304})+$signed(-{1'b0,x249})+$signed(-{1'b0,x121});
assign sharing50 = $signed(-{1'b0,x229})+$signed(-{1'b0,x237})+$signed({1'b0,x228})+$signed(-{1'b0,x108})+$signed(-{1'b0,x292})+$signed(-{1'b0,x109});
assign sharing51 = $signed(-{1'b0,x110})+$signed(-{1'b0,x231})+$signed(-{1'b0,x239})+$signed({1'b0,x230})+$signed(-{1'b0,x294})+$signed(-{1'b0,x111});
assign sharing52 = $signed(-{1'b0,x126})+$signed(-{1'b0,x255})+$signed(-{1'b0,x247})+$signed({1'b0,x246})+$signed(-{1'b0,x310})+$signed(-{1'b0,x127});
assign sharing53 = $signed(-{1'b0,x106})+$signed(-{1'b0,x227})+$signed(-{1'b0,x107})+$signed({1'b0,x226})+$signed(-{1'b0,x290})+$signed(-{1'b0,x235});
assign sharing54 = $signed({1'b0,x192})+$signed(-{1'b0,x72})+$signed(-{1'b0,x256})+$signed(-{1'b0,x73})+$signed(-{1'b0,x193})+$signed(-{1'b0,x201});
assign sharing55 = $signed(-{1'b0,x90})+$signed(-{1'b0,x211})+$signed(-{1'b0,x219})+$signed(-{1'b0,x274})+$signed({1'b0,x210})+$signed(-{1'b0,x91});
assign sharing56 = $signed(-{1'b0,x78})+$signed(-{1'b0,x199})+$signed(-{1'b0,x207})+$signed(-{1'b0,x262})+$signed({1'b0,x198})+$signed(-{1'b0,x79});
assign sharing57 = $signed(-{1'b0,x94})+$signed(-{1'b0,x215})+$signed(-{1'b0,x223})+$signed(-{1'b0,x278})+$signed({1'b0,x214})+$signed(-{1'b0,x95});
assign sharing58 = $signed(-{1'b0,x225})+$signed(-{1'b0,x105})+$signed({1'b0,x224})+$signed(-{1'b0,x104})+$signed(-{1'b0,x288})+$signed(-{1'b0,x233});
assign sharing59 = $signed(-{1'b0,x122})+$signed(-{1'b0,x251})+$signed(-{1'b0,x243})+$signed({1'b0,x242})+$signed(-{1'b0,x306})+$signed(-{1'b0,x123});
assign sharing60 = $signed(-{1'b0,x74})+$signed(-{1'b0,x195})+$signed(-{1'b0,x203})+$signed(-{1'b0,x258})+$signed({1'b0,x194})+$signed(-{1'b0,x75});
assign sharing61 = $signed({1'b0,x212})+$signed(-{1'b0,x92})+$signed(-{1'b0,x276})+$signed(-{1'b0,x213})+$signed(-{1'b0,x93})+$signed(-{1'b0,x221});
assign sharing62 = $signed({1'b0,x208})+$signed(-{1'b0,x88})+$signed(-{1'b0,x272})+$signed(-{1'b0,x89})+$signed(-{1'b0,x209})+$signed(-{1'b0,x217});
assign sharing63 = $signed({1'b0,x196})+$signed(-{1'b0,x76})+$signed(-{1'b0,x260})+$signed(-{1'b0,x205})+$signed(-{1'b0,x197})+$signed(-{1'b0,x77});
assign sharing64 = $signed(-{1'b0,x245})+$signed({1'b0,x244})+$signed(-{1'b0,x124})+$signed(-{1'b0,x308})+$signed(-{1'b0,x253})+$signed(-{1'b0,x125});
assign sharing65 = $signed(-{1'b0,x36})+$signed(-{2'b0,x165}<<<3'd1)+$signed({1'b0,x45});
assign sharing66 = $signed(-{1'b0,x365})+$signed(-{2'b0,x300}<<<3'd1)+$signed(-{2'b0,x364}<<<3'd1)+$signed({2'b0,x173}<<<3'd1)+$signed({2'b0,x293}<<<3'd1)+$signed(-{1'b0,x37});
assign sharing67 = $signed(-{2'b0,x64}<<<3'd1)+$signed(-{1'b0,x264})+$signed(-{1'b0,x320})+$signed({1'b0,x137})+$signed(-{2'b0,x72}<<<3'd1)+$signed({1'b0,x129})+$signed(-{2'b0,x65}<<<3'd1);
assign sharing68 = $signed(-{1'b0,x6})+$signed(-{2'b0,x135}<<<3'd1)+$signed({1'b0,x15});
assign sharing69 = $signed(-{1'b0,x335})+$signed({2'b0,x263}<<<3'd1)+$signed(-{2'b0,x270}<<<3'd1)+$signed(-{2'b0,x334}<<<3'd1)+$signed({2'b0,x143}<<<3'd1)+$signed(-{1'b0,x7});
assign sharing70 = $signed(-{1'b0,x32})+$signed(-{2'b0,x161}<<<3'd1)+$signed({1'b0,x41});
assign sharing71 = $signed(-{1'b0,x361})+$signed(-{2'b0,x296}<<<3'd1)+$signed(-{2'b0,x360}<<<3'd1)+$signed({2'b0,x169}<<<3'd1)+$signed({2'b0,x289}<<<3'd1)+$signed(-{1'b0,x33});
assign sharing72 = $signed(-{1'b0,x2})+$signed(-{2'b0,x131}<<<3'd1)+$signed({1'b0,x11});
assign sharing73 = $signed(-{1'b0,x331})+$signed({2'b0,x259}<<<3'd1)+$signed(-{2'b0,x266}<<<3'd1)+$signed(-{2'b0,x330}<<<3'd1)+$signed({2'b0,x139}<<<3'd1)+$signed(-{1'b0,x3});
assign sharing74 = $signed(-{1'b0,x20})+$signed(-{2'b0,x149}<<<3'd1)+$signed({1'b0,x29});
assign sharing75 = $signed(-{2'b0,x284}<<<3'd1)+$signed(-{2'b0,x348}<<<3'd1)+$signed({2'b0,x157}<<<3'd1)+$signed({2'b0,x277}<<<3'd1)+$signed(-{1'b0,x21})+$signed(-{1'b0,x349});
assign sharing76 = $signed(-{1'b0,x16})+$signed(-{2'b0,x145}<<<3'd1)+$signed({1'b0,x25});
assign sharing77 = $signed({2'b0,x280}<<<3'd1)+$signed({2'b0,x344}<<<3'd1)+$signed(-{2'b0,x153}<<<3'd1)+$signed({1'b0,x17})+$signed(-{2'b0,x273}<<<3'd1)+$signed({1'b0,x345});
assign sharing78 = $signed({2'b0,x80}<<<3'd1)+$signed({1'b0,x280})+$signed({1'b0,x336})+$signed({2'b0,x88}<<<3'd1)+$signed({2'b0,x81}<<<3'd1)+$signed(-{1'b0,x145})+$signed(-{1'b0,x153});
assign sharing79 = $signed({2'b0,x68}<<<3'd1)+$signed({1'b0,x268})+$signed({1'b0,x324})+$signed({2'b0,x76}<<<3'd1)+$signed({2'b0,x69}<<<3'd1)+$signed(-{1'b0,x133})+$signed(-{1'b0,x141});
assign sharing80 = $signed({2'b0,x114}<<<3'd1)+$signed(-{1'b0,x179})+$signed(-{1'b0,x187})+$signed({2'b0,x122}<<<3'd1)+$signed({1'b0,x370})+$signed({2'b0,x115}<<<3'd1)+$signed({1'b0,x314});
assign sharing81 = $signed(-{1'b0,x48})+$signed(-{2'b0,x177}<<<3'd1)+$signed({1'b0,x57});
assign sharing82 = $signed({2'b0,x312}<<<3'd1)+$signed({2'b0,x376}<<<3'd1)+$signed({1'b0,x377})+$signed(-{2'b0,x305}<<<3'd1)+$signed({1'b0,x49})+$signed(-{2'b0,x185}<<<3'd1);
assign sharing83 = $signed(-{2'b0,x104}<<<3'd1)+$signed(-{1'b0,x296})+$signed(-{1'b0,x352})+$signed(-{2'b0,x96}<<<3'd1)+$signed(-{2'b0,x97}<<<3'd1)+$signed({1'b0,x161})+$signed({1'b0,x169});
assign sharing84 = $signed(-{1'b0,x38})+$signed(-{2'b0,x167}<<<3'd1)+$signed({1'b0,x47});
assign sharing85 = $signed(-{2'b0,x366}<<<3'd1)+$signed(-{1'b0,x367})+$signed(-{2'b0,x302}<<<3'd1)+$signed({2'b0,x295}<<<3'd1)+$signed({2'b0,x175}<<<3'd1)+$signed(-{1'b0,x39});
assign sharing86 = $signed(-{2'b0,x84}<<<3'd1)+$signed(-{1'b0,x284})+$signed({1'b0,x157})+$signed(-{1'b0,x340})+$signed(-{2'b0,x92}<<<3'd1)+$signed({1'b0,x149})+$signed(-{2'b0,x85}<<<3'd1);
assign sharing87 = $signed(-{1'b0,x34})+$signed(-{2'b0,x163}<<<3'd1)+$signed({1'b0,x43});
assign sharing88 = $signed(-{2'b0,x362}<<<3'd1)+$signed(-{1'b0,x363})+$signed(-{2'b0,x298}<<<3'd1)+$signed({2'b0,x291}<<<3'd1)+$signed({2'b0,x171}<<<3'd1)+$signed(-{1'b0,x35});
assign sharing89 = $signed(-{1'b0,x52})+$signed(-{2'b0,x181}<<<3'd1)+$signed({1'b0,x61});
assign sharing90 = $signed(-{2'b0,x316}<<<3'd1)+$signed(-{2'b0,x380}<<<3'd1)+$signed(-{1'b0,x381})+$signed({2'b0,x309}<<<3'd1)+$signed({2'b0,x189}<<<3'd1)+$signed(-{1'b0,x53});
assign sharing91 = $signed({2'b0,x87}<<<3'd1)+$signed({1'b0,x286})+$signed({2'b0,x86}<<<3'd1)+$signed({1'b0,x342})+$signed(-{1'b0,x159})+$signed({2'b0,x94}<<<3'd1)+$signed(-{1'b0,x151});
assign sharing92 = $signed(-{1'b0,x4})+$signed(-{2'b0,x133}<<<3'd1)+$signed({1'b0,x13});
assign sharing93 = $signed(-{2'b0,x268}<<<3'd1)+$signed(-{2'b0,x332}<<<3'd1)+$signed(-{1'b0,x5})+$signed({2'b0,x141}<<<3'd1)+$signed({2'b0,x261}<<<3'd1)+$signed(-{1'b0,x333});
assign sharing94 = $signed(-{1'b0,x22})+$signed(-{2'b0,x151}<<<3'd1)+$signed({1'b0,x31});
assign sharing95 = $signed(-{1'b0,x351})+$signed(-{2'b0,x350}<<<3'd1)+$signed({2'b0,x279}<<<3'd1)+$signed(-{2'b0,x286}<<<3'd1)+$signed({2'b0,x159}<<<3'd1)+$signed(-{1'b0,x23});
assign sharing96 = $signed(-{1'b0,x326})+$signed(-{2'b0,x70}<<<3'd1)+$signed(-{2'b0,x78}<<<3'd1)+$signed(-{1'b0,x270})+$signed({1'b0,x143})+$signed(-{2'b0,x71}<<<3'd1)+$signed({1'b0,x135});
assign sharing97 = $signed(-{1'b0,x0})+$signed(-{2'b0,x129}<<<3'd1)+$signed({1'b0,x9});
assign sharing98 = $signed(-{2'b0,x264}<<<3'd1)+$signed(-{2'b0,x328}<<<3'd1)+$signed(-{1'b0,x1})+$signed({2'b0,x137}<<<3'd1)+$signed({2'b0,x257}<<<3'd1)+$signed(-{1'b0,x329});
assign sharing99 = $signed({2'b0,x120}<<<3'd1)+$signed({2'b0,x112}<<<3'd1)+$signed({1'b0,x368})+$signed({1'b0,x312})+$signed({2'b0,x113}<<<3'd1)+$signed(-{1'b0,x177})+$signed(-{1'b0,x185});
assign sharing100 = $signed({2'b0,x83}<<<3'd1)+$signed({1'b0,x338})+$signed({2'b0,x82}<<<3'd1)+$signed({1'b0,x282})+$signed(-{1'b0,x155})+$signed({2'b0,x90}<<<3'd1)+$signed(-{1'b0,x147});
assign sharing101 = $signed(-{1'b0,x18})+$signed(-{2'b0,x147}<<<3'd1)+$signed({1'b0,x27});
assign sharing102 = $signed(-{1'b0,x347})+$signed(-{2'b0,x346}<<<3'd1)+$signed({2'b0,x275}<<<3'd1)+$signed(-{2'b0,x282}<<<3'd1)+$signed({2'b0,x155}<<<3'd1)+$signed(-{1'b0,x19});
assign sharing103 = $signed(-{1'b0,x322})+$signed(-{2'b0,x66}<<<3'd1)+$signed(-{1'b0,x266})+$signed(-{2'b0,x74}<<<3'd1)+$signed({1'b0,x139})+$signed(-{2'b0,x67}<<<3'd1)+$signed({1'b0,x131});
assign sharing104 = $signed({2'b0,x108}<<<3'd1)+$signed({1'b0,x300})+$signed({1'b0,x356})+$signed({2'b0,x100}<<<3'd1)+$signed({2'b0,x101}<<<3'd1)+$signed(-{1'b0,x165})+$signed(-{1'b0,x173});
assign sharing105 = $signed({2'b0,x118}<<<3'd1)+$signed(-{1'b0,x183})+$signed(-{1'b0,x191})+$signed({2'b0,x126}<<<3'd1)+$signed({1'b0,x374})+$signed({2'b0,x119}<<<3'd1)+$signed({1'b0,x318});
assign sharing106 = $signed(-{1'b0,x54})+$signed(-{2'b0,x183}<<<3'd1)+$signed({1'b0,x63});
assign sharing107 = $signed(-{2'b0,x382}<<<3'd1)+$signed({2'b0,x191}<<<3'd1)+$signed(-{2'b0,x318}<<<3'd1)+$signed(-{1'b0,x383})+$signed({2'b0,x311}<<<3'd1)+$signed(-{1'b0,x55});
assign sharing108 = $signed(-{2'b0,x110}<<<3'd1)+$signed({1'b0,x175})+$signed(-{1'b0,x358})+$signed(-{2'b0,x102}<<<3'd1)+$signed(-{1'b0,x302})+$signed(-{2'b0,x103}<<<3'd1)+$signed({1'b0,x167});
assign sharing109 = $signed(-{1'b0,x50})+$signed(-{2'b0,x179}<<<3'd1)+$signed({1'b0,x59});
assign sharing110 = $signed(-{2'b0,x378}<<<3'd1)+$signed({2'b0,x187}<<<3'd1)+$signed(-{2'b0,x314}<<<3'd1)+$signed(-{1'b0,x379})+$signed({2'b0,x307}<<<3'd1)+$signed(-{1'b0,x51});
assign sharing111 = $signed({1'b0,x171})+$signed(-{1'b0,x354})+$signed(-{2'b0,x106}<<<3'd1)+$signed(-{1'b0,x298})+$signed(-{2'b0,x98}<<<3'd1)+$signed(-{2'b0,x99}<<<3'd1)+$signed({1'b0,x163});
assign sharing112 = $signed(-{2'b0,x124}<<<3'd1)+$signed(-{2'b0,x116}<<<3'd1)+$signed(-{1'b0,x372})+$signed(-{1'b0,x316})+$signed(-{2'b0,x117}<<<3'd1)+$signed({1'b0,x181})+$signed({1'b0,x189});
wire signed[11:0] temp_y  [0:207];
assign temp_y[0] = 
$signed(-{3'b0,x328}<<<3'd2)+$signed({2'b0,x264}<<<3'd1)+$signed(-{2'b0,x320}<<<3'd1)+$signed(-{1'b0,x72})+$signed({1'b0,x136})+$signed({2'b0,x257}<<<3'd1)+$signed({1'b0,x265})+$signed(-{1'b0,x73})+$signed(-{1'b0,x129})+$signed(-{3'b0,x329}<<<3'd2)+$signed(sharing45)+$signed(11'd32);
assign y0=temp_y[0][11] ==1'b1 ? 5'd0 :  
        temp_y[0][9] ==1'b1 ? 5'd31 : 
        temp_y[0][3]==1'b1 ? temp_y[0][8:4]+1'b1 : temp_y[0][8:4];
assign temp_y[1] = 
$signed({2'b0,x72}<<<3'd1)+$signed({1'b0,x0})+$signed({1'b0,x64})+$signed({2'b0,x200}<<<3'd1)+$signed({2'b0,x328}<<<3'd1)+$signed(-{1'b0,x264})+$signed(-{1'b0,x1})+$signed(-{2'b0,x201}<<<3'd1)+$signed(-{1'b0,x257})+$signed(-{1'b0,x136})+$signed({3'b0,x329}<<<3'd2)+$signed(sharing45)-$signed(11'd0);
assign y1=temp_y[1][11] ==1'b1 ? 5'd0 :  
        temp_y[1][9] ==1'b1 ? 5'd31 : 
        temp_y[1][3]==1'b1 ? temp_y[1][8:4]+1'b1 : temp_y[1][8:4];
assign temp_y[2] = 
$signed(-{3'b0,x256}<<<3'd2)+$signed(-{2'b0,x64}<<<3'd1)+$signed({1'b0,x128})+$signed(-{2'b0,x72}<<<3'd1)+$signed(-{4'b0,x257}<<<3'd3)+$signed(-{3'b0,x264}<<<3'd2)+$signed(-{3'b0,x265}<<<3'd2)+$signed(-{2'b0,x320}<<<3'd1)+$signed(sharing21)+$signed(sharing22)+$signed(11'd40);
assign y2=temp_y[2][11] ==1'b1 ? 5'd0 :  
        temp_y[2][9] ==1'b1 ? 5'd31 : 
        temp_y[2][3]==1'b1 ? temp_y[2][8:4]+1'b1 : temp_y[2][8:4];
assign temp_y[3] = 
$signed({2'b0,x320}<<<3'd1)+$signed({1'b0,x256})+$signed({1'b0,x8})+$signed({1'b0,x136})+$signed(-{1'b0,x64})+$signed({1'b0,x265})+$signed({1'b0,x321})+$signed(-{1'b0,x192})+$signed(-{1'b0,x72})+$signed(-{2'b0,x73}<<<3'd1)+$signed(sharing97)+$signed(sharing98)-$signed(11'd16);
assign y3=temp_y[3][11] ==1'b1 ? 5'd0 :  
        temp_y[3][9] ==1'b1 ? 5'd31 : 
        temp_y[3][3]==1'b1 ? temp_y[3][8:4]+1'b1 : temp_y[3][8:4];
assign temp_y[4] = 
$signed({3'b0,x136}<<<3'd2)+$signed(-{2'b0,x128}<<<3'd1)+$signed({1'b0,x320})+$signed(-{2'b0,x8}<<<3'd1)+$signed(-{1'b0,x200})+$signed(-{2'b0,x201}<<<3'd1)+$signed(-{2'b0,x65}<<<3'd1)+$signed(-{2'b0,x321}<<<3'd1)+$signed(sharing97)+$signed(-sharing98)-$signed(11'd24);
assign y4=temp_y[4][11] ==1'b1 ? 5'd0 :  
        temp_y[4][9] ==1'b1 ? 5'd31 : 
        temp_y[4][3]==1'b1 ? temp_y[4][8:4]+1'b1 : temp_y[4][8:4];
assign temp_y[5] = 
$signed({2'b0,x256}<<<3'd1)+$signed({1'b0,x200})+$signed({2'b0,x128}<<<3'd1)+$signed({2'b0,x264}<<<3'd1)+$signed({3'b0,x265}<<<3'd2)+$signed({1'b0,x201})+$signed(-{1'b0,x192})+$signed(-{1'b0,x72})+$signed(-{1'b0,x0})+$signed(-{1'b0,x320})+$signed(-{1'b0,x193})+$signed(-{1'b0,x1})+$signed(-{1'b0,x329})-$signed(11'd32);
assign y5=temp_y[5][11] ==1'b1 ? 5'd0 :  
        temp_y[5][9] ==1'b1 ? 5'd31 : 
        temp_y[5][3]==1'b1 ? temp_y[5][8:4]+1'b1 : temp_y[5][8:4];
assign temp_y[6] = 
$signed(-{1'b0,x64})+$signed({3'b0,x321}<<<3'd2)+$signed(-{2'b0,x265}<<<3'd1)+$signed({3'b0,x329}<<<3'd2)+$signed(-{2'b0,x257}<<<3'd1)+$signed(-{1'b0,x1})+$signed(-{1'b0,x9})+$signed(sharing54)-$signed(11'd0);
assign y6=temp_y[6][11] ==1'b1 ? 5'd0 :  
        temp_y[6][9] ==1'b1 ? 5'd31 : 
        temp_y[6][3]==1'b1 ? temp_y[6][8:4]+1'b1 : temp_y[6][8:4];
assign temp_y[7] = 
$signed(-{2'b0,x256}<<<3'd1)+$signed(-{1'b0,x128})+$signed({1'b0,x192})+$signed({3'b0,x73}<<<3'd2)+$signed({2'b0,x321}<<<3'd1)+$signed({1'b0,x257})+$signed(-{3'b0,x329}<<<3'd2)+$signed(-{1'b0,x193})+$signed(-{1'b0,x328})+$signed(-sharing67)-$signed(11'd0);
assign y7=temp_y[7][11] ==1'b1 ? 5'd0 :  
        temp_y[7][9] ==1'b1 ? 5'd31 : 
        temp_y[7][3]==1'b1 ? temp_y[7][8:4]+1'b1 : temp_y[7][8:4];
assign temp_y[8] = 
$signed(-{3'b0,x8}<<<3'd2)+$signed(-{2'b0,x192}<<<3'd1)+$signed({1'b0,x328})+$signed(-{1'b0,x136})+$signed(-{1'b0,x264})+$signed({2'b0,x193}<<<3'd1)+$signed(-{2'b0,x9}<<<3'd1)+$signed(-{2'b0,x137}<<<3'd1)+$signed(-{2'b0,x0}<<<3'd1)+$signed({1'b0,x64})+$signed(sharing2)+$signed(11'd40);
assign y8=temp_y[8][11] ==1'b1 ? 5'd0 :  
        temp_y[8][9] ==1'b1 ? 5'd31 : 
        temp_y[8][3]==1'b1 ? temp_y[8][8:4]+1'b1 : temp_y[8][8:4];
assign temp_y[9] = 
$signed(-{2'b0,x8}<<<3'd1)+$signed({1'b0,x192})+$signed({4'b0,x9}<<<3'd3)+$signed(-{2'b0,x0}<<<3'd1)+$signed(-{2'b0,x201}<<<3'd1)+$signed(-{1'b0,x329})+$signed(-{1'b0,x193})+$signed({1'b0,x64})+$signed(-sharing2)-$signed(11'd8);
assign y9=temp_y[9][11] ==1'b1 ? 5'd0 :  
        temp_y[9][9] ==1'b1 ? 5'd31 : 
        temp_y[9][3]==1'b1 ? temp_y[9][8:4]+1'b1 : temp_y[9][8:4];
assign temp_y[10] = 
$signed({3'b0,x320}<<<3'd2)+$signed(-{2'b0,x128}<<<3'd1)+$signed(-{2'b0,x0}<<<3'd1)+$signed(-{1'b0,x72})+$signed(-{1'b0,x8})+$signed({2'b0,x9}<<<3'd1)+$signed({2'b0,x129}<<<3'd1)+$signed(-{1'b0,x136})+$signed(-{1'b0,x73})+$signed(-{1'b0,x65})+$signed(-{2'b0,x256}<<<3'd1)+$signed(-{1'b0,x257})+$signed(-{2'b0,x265}<<<3'd1)+$signed(-{1'b0,x264})+$signed(sharing21)+$signed(-sharing22)-$signed(11'd16);
assign y10=temp_y[10][11] ==1'b1 ? 5'd0 :  
        temp_y[10][9] ==1'b1 ? 5'd31 : 
        temp_y[10][3]==1'b1 ? temp_y[10][8:4]+1'b1 : temp_y[10][8:4];
assign temp_y[11] = 
$signed(-{4'b0,x264}<<<3'd3)+$signed(-{3'b0,x192}<<<3'd2)+$signed(-{3'b0,x256}<<<3'd2)+$signed(-{1'b0,x200})+$signed(-{4'b0,x257}<<<3'd3)+$signed(-{4'b0,x201}<<<3'd3)+$signed(-{1'b0,x319})+$signed({1'b0,x9})+$signed(-{1'b0,x73})+$signed(-{1'b0,x193})+$signed(-{1'b0,x328})+$signed(-{1'b0,x327})+$signed(sharing67)+$signed(11'd24);
assign y11=temp_y[11][11] ==1'b1 ? 5'd0 :  
        temp_y[11][9] ==1'b1 ? 5'd31 : 
        temp_y[11][3]==1'b1 ? temp_y[11][8:4]+1'b1 : temp_y[11][8:4];
assign temp_y[12] = 
$signed({3'b0,x200}<<<3'd2)+$signed({2'b0,x128}<<<3'd1)+$signed({2'b0,x320}<<<3'd1)+$signed(-{2'b0,x264}<<<3'd1)+$signed({1'b0,x328})+$signed(-{1'b0,x8})+$signed(-{1'b0,x257})+$signed(-{3'b0,x137}<<<3'd2)+$signed(-{3'b0,x129}<<<3'd2)+$signed(-{2'b0,x65}<<<3'd1)+$signed(-{1'b0,x321})+$signed({1'b0,x9})+$signed({1'b0,x64})+$signed(sharing54)+$signed(11'd16);
assign y12=temp_y[12][11] ==1'b1 ? 5'd0 :  
        temp_y[12][9] ==1'b1 ? 5'd31 : 
        temp_y[12][3]==1'b1 ? temp_y[12][8:4]+1'b1 : temp_y[12][8:4];
assign temp_y[13] = 
$signed(-{3'b0,x330}<<<3'd2)+$signed({2'b0,x266}<<<3'd1)+$signed(-{2'b0,x322}<<<3'd1)+$signed(-{1'b0,x74})+$signed({1'b0,x138})+$signed({2'b0,x259}<<<3'd1)+$signed({1'b0,x267})+$signed(-{1'b0,x75})+$signed(-{1'b0,x131})+$signed(-{3'b0,x331}<<<3'd2)+$signed(sharing37)+$signed(11'd32);
assign y13=temp_y[13][11] ==1'b1 ? 5'd0 :  
        temp_y[13][9] ==1'b1 ? 5'd31 : 
        temp_y[13][3]==1'b1 ? temp_y[13][8:4]+1'b1 : temp_y[13][8:4];
assign temp_y[14] = 
$signed({2'b0,x74}<<<3'd1)+$signed({1'b0,x66})+$signed({1'b0,x2})+$signed({2'b0,x202}<<<3'd1)+$signed({2'b0,x330}<<<3'd1)+$signed(-{1'b0,x266})+$signed(-{1'b0,x3})+$signed(-{2'b0,x203}<<<3'd1)+$signed(-{1'b0,x259})+$signed(-{1'b0,x138})+$signed({3'b0,x331}<<<3'd2)+$signed(sharing37)-$signed(11'd0);
assign y14=temp_y[14][11] ==1'b1 ? 5'd0 :  
        temp_y[14][9] ==1'b1 ? 5'd31 : 
        temp_y[14][3]==1'b1 ? temp_y[14][8:4]+1'b1 : temp_y[14][8:4];
assign temp_y[15] = 
$signed(-{3'b0,x258}<<<3'd2)+$signed({2'b0,x202}<<<3'd1)+$signed({1'b0,x130})+$signed({1'b0,x194})+$signed(-{2'b0,x66}<<<3'd1)+$signed(-{2'b0,x74}<<<3'd1)+$signed(-{4'b0,x259}<<<3'd3)+$signed(-{3'b0,x266}<<<3'd2)+$signed(-{3'b0,x267}<<<3'd2)+$signed(-{1'b0,x203})+$signed(-{1'b0,x139})+$signed(-{3'b0,x330}<<<3'd2)+$signed(-{2'b0,x322}<<<3'd1)+$signed(11'd40);
assign y15=temp_y[15][11] ==1'b1 ? 5'd0 :  
        temp_y[15][9] ==1'b1 ? 5'd31 : 
        temp_y[15][3]==1'b1 ? temp_y[15][8:4]+1'b1 : temp_y[15][8:4];
assign temp_y[16] = 
$signed({2'b0,x322}<<<3'd1)+$signed(-{1'b0,x66})+$signed({1'b0,x10})+$signed({1'b0,x258})+$signed({1'b0,x138})+$signed({1'b0,x323})+$signed({1'b0,x267})+$signed(-{1'b0,x194})+$signed(-{1'b0,x74})+$signed(-{2'b0,x75}<<<3'd1)+$signed(sharing72)+$signed(sharing73)-$signed(11'd16);
assign y16=temp_y[16][11] ==1'b1 ? 5'd0 :  
        temp_y[16][9] ==1'b1 ? 5'd31 : 
        temp_y[16][3]==1'b1 ? temp_y[16][8:4]+1'b1 : temp_y[16][8:4];
assign temp_y[17] = 
$signed({3'b0,x138}<<<3'd2)+$signed(-{2'b0,x130}<<<3'd1)+$signed({1'b0,x322})+$signed(-{2'b0,x10}<<<3'd1)+$signed(-{1'b0,x202})+$signed(-{2'b0,x203}<<<3'd1)+$signed(-{2'b0,x67}<<<3'd1)+$signed(-{2'b0,x323}<<<3'd1)+$signed(sharing72)+$signed(-sharing73)-$signed(11'd24);
assign y17=temp_y[17][11] ==1'b1 ? 5'd0 :  
        temp_y[17][9] ==1'b1 ? 5'd31 : 
        temp_y[17][3]==1'b1 ? temp_y[17][8:4]+1'b1 : temp_y[17][8:4];
assign temp_y[18] = 
$signed({2'b0,x266}<<<3'd1)+$signed(-{1'b0,x2})+$signed(-{1'b0,x322})+$signed({1'b0,x202})+$signed({3'b0,x267}<<<3'd2)+$signed(-{1'b0,x195})+$signed(-{1'b0,x331})+$signed(-{1'b0,x3})+$signed(-{1'b0,x74})+$signed(-{1'b0,x194})+$signed(sharing12)-$signed(11'd32);
assign y18=temp_y[18][11] ==1'b1 ? 5'd0 :  
        temp_y[18][9] ==1'b1 ? 5'd31 : 
        temp_y[18][3]==1'b1 ? temp_y[18][8:4]+1'b1 : temp_y[18][8:4];
assign temp_y[19] = 
$signed(-{1'b0,x66})+$signed({3'b0,x331}<<<3'd2)+$signed({3'b0,x323}<<<3'd2)+$signed(-{1'b0,x3})+$signed(-{2'b0,x267}<<<3'd1)+$signed(-{2'b0,x259}<<<3'd1)+$signed(-{1'b0,x11})+$signed(sharing60)-$signed(11'd0);
assign y19=temp_y[19][11] ==1'b1 ? 5'd0 :  
        temp_y[19][9] ==1'b1 ? 5'd31 : 
        temp_y[19][3]==1'b1 ? temp_y[19][8:4]+1'b1 : temp_y[19][8:4];
assign temp_y[20] = 
$signed(-{2'b0,x258}<<<3'd1)+$signed({1'b0,x194})+$signed(-{1'b0,x130})+$signed({3'b0,x75}<<<3'd2)+$signed(-{3'b0,x331}<<<3'd2)+$signed({2'b0,x323}<<<3'd1)+$signed({1'b0,x259})+$signed(-{1'b0,x195})+$signed(-{1'b0,x330})+$signed(-sharing103)-$signed(11'd0);
assign y20=temp_y[20][11] ==1'b1 ? 5'd0 :  
        temp_y[20][9] ==1'b1 ? 5'd31 : 
        temp_y[20][3]==1'b1 ? temp_y[20][8:4]+1'b1 : temp_y[20][8:4];
assign temp_y[21] = 
$signed(-{3'b0,x10}<<<3'd2)+$signed(-{2'b0,x194}<<<3'd1)+$signed({1'b0,x330})+$signed(-{1'b0,x138})+$signed(-{1'b0,x266})+$signed({2'b0,x195}<<<3'd1)+$signed(-{2'b0,x11}<<<3'd1)+$signed(-{2'b0,x139}<<<3'd1)+$signed(-{2'b0,x2}<<<3'd1)+$signed({1'b0,x66})+$signed(sharing16)+$signed(11'd40);
assign y21=temp_y[21][11] ==1'b1 ? 5'd0 :  
        temp_y[21][9] ==1'b1 ? 5'd31 : 
        temp_y[21][3]==1'b1 ? temp_y[21][8:4]+1'b1 : temp_y[21][8:4];
assign temp_y[22] = 
$signed(-{2'b0,x10}<<<3'd1)+$signed({1'b0,x194})+$signed({4'b0,x11}<<<3'd3)+$signed(-{2'b0,x2}<<<3'd1)+$signed(-{2'b0,x203}<<<3'd1)+$signed(-{1'b0,x195})+$signed(-{1'b0,x331})+$signed({1'b0,x66})+$signed(-sharing16)-$signed(11'd8);
assign y22=temp_y[22][11] ==1'b1 ? 5'd0 :  
        temp_y[22][9] ==1'b1 ? 5'd31 : 
        temp_y[22][3]==1'b1 ? temp_y[22][8:4]+1'b1 : temp_y[22][8:4];
assign temp_y[23] = 
$signed(-{1'b0,x74})+$signed({3'b0,x330}<<<3'd2)+$signed(-{2'b0,x2}<<<3'd1)+$signed(-{1'b0,x138})+$signed({3'b0,x322}<<<3'd2)+$signed(-{1'b0,x10})+$signed({2'b0,x11}<<<3'd1)+$signed({2'b0,x131}<<<3'd1)+$signed({1'b0,x139})+$signed(-{2'b0,x202}<<<3'd1)+$signed(-{2'b0,x267}<<<3'd1)+$signed(-{1'b0,x67})+$signed(-{1'b0,x75})+$signed(-{1'b0,x259})+$signed(-{1'b0,x194})+$signed(-{1'b0,x266})+$signed(-sharing12)-$signed(11'd16);
assign y23=temp_y[23][11] ==1'b1 ? 5'd0 :  
        temp_y[23][9] ==1'b1 ? 5'd31 : 
        temp_y[23][3]==1'b1 ? temp_y[23][8:4]+1'b1 : temp_y[23][8:4];
assign temp_y[24] = 
$signed(-{1'b0,x321})+$signed(-{4'b0,x266}<<<3'd3)+$signed(-{3'b0,x194}<<<3'd2)+$signed(-{3'b0,x258}<<<3'd2)+$signed(-{1'b0,x329})+$signed(-{4'b0,x259}<<<3'd3)+$signed(-{1'b0,x202})+$signed(-{4'b0,x203}<<<3'd3)+$signed({1'b0,x11})+$signed(-{1'b0,x75})+$signed(-{1'b0,x195})+$signed(-{1'b0,x330})+$signed(sharing103)+$signed(11'd24);
assign y24=temp_y[24][11] ==1'b1 ? 5'd0 :  
        temp_y[24][9] ==1'b1 ? 5'd31 : 
        temp_y[24][3]==1'b1 ? temp_y[24][8:4]+1'b1 : temp_y[24][8:4];
assign temp_y[25] = 
$signed({1'b0,x66})+$signed({3'b0,x202}<<<3'd2)+$signed({2'b0,x130}<<<3'd1)+$signed({2'b0,x322}<<<3'd1)+$signed({1'b0,x330})+$signed(-{3'b0,x131}<<<3'd2)+$signed(-{2'b0,x266}<<<3'd1)+$signed(-{1'b0,x323})+$signed(-{1'b0,x10})+$signed(-{3'b0,x139}<<<3'd2)+$signed(-{2'b0,x67}<<<3'd1)+$signed(-{1'b0,x259})+$signed({1'b0,x11})+$signed(sharing60)+$signed(11'd16);
assign y25=temp_y[25][11] ==1'b1 ? 5'd0 :  
        temp_y[25][9] ==1'b1 ? 5'd31 : 
        temp_y[25][3]==1'b1 ? temp_y[25][8:4]+1'b1 : temp_y[25][8:4];
assign temp_y[26] = 
$signed(-{3'b0,x332}<<<3'd2)+$signed({2'b0,x268}<<<3'd1)+$signed(-{2'b0,x324}<<<3'd1)+$signed(-{1'b0,x76})+$signed({1'b0,x269})+$signed({2'b0,x261}<<<3'd1)+$signed(-{1'b0,x133})+$signed({1'b0,x140})+$signed(-{3'b0,x333}<<<3'd2)+$signed(-{1'b0,x77})+$signed(sharing40)+$signed(11'd32);
assign y26=temp_y[26][11] ==1'b1 ? 5'd0 :  
        temp_y[26][9] ==1'b1 ? 5'd31 : 
        temp_y[26][3]==1'b1 ? temp_y[26][8:4]+1'b1 : temp_y[26][8:4];
assign temp_y[27] = 
$signed({2'b0,x76}<<<3'd1)+$signed({1'b0,x4})+$signed({1'b0,x68})+$signed({2'b0,x204}<<<3'd1)+$signed({2'b0,x332}<<<3'd1)+$signed(-{1'b0,x268})+$signed(-{1'b0,x261})+$signed(-{2'b0,x205}<<<3'd1)+$signed(-{1'b0,x5})+$signed(-{1'b0,x140})+$signed({3'b0,x333}<<<3'd2)+$signed(sharing40)-$signed(11'd0);
assign y27=temp_y[27][11] ==1'b1 ? 5'd0 :  
        temp_y[27][9] ==1'b1 ? 5'd31 : 
        temp_y[27][3]==1'b1 ? temp_y[27][8:4]+1'b1 : temp_y[27][8:4];
assign temp_y[28] = 
$signed(-{1'b0,x141})+$signed(-{3'b0,x260}<<<3'd2)+$signed({2'b0,x204}<<<3'd1)+$signed({1'b0,x132})+$signed({1'b0,x196})+$signed(-{2'b0,x68}<<<3'd1)+$signed(-{2'b0,x76}<<<3'd1)+$signed(-{1'b0,x205})+$signed(-{4'b0,x261}<<<3'd3)+$signed(-{3'b0,x268}<<<3'd2)+$signed(-{3'b0,x269}<<<3'd2)+$signed(-{2'b0,x324}<<<3'd1)+$signed(-{3'b0,x332}<<<3'd2)+$signed(11'd40);
assign y28=temp_y[28][11] ==1'b1 ? 5'd0 :  
        temp_y[28][9] ==1'b1 ? 5'd31 : 
        temp_y[28][3]==1'b1 ? temp_y[28][8:4]+1'b1 : temp_y[28][8:4];
assign temp_y[29] = 
$signed({2'b0,x324}<<<3'd1)+$signed({1'b0,x260})+$signed({1'b0,x12})+$signed({1'b0,x140})+$signed(-{1'b0,x68})+$signed({1'b0,x269})+$signed(-{1'b0,x196})+$signed(-{1'b0,x76})+$signed(-{2'b0,x77}<<<3'd1)+$signed({1'b0,x325})+$signed(sharing92)+$signed(sharing93)-$signed(11'd16);
assign y29=temp_y[29][11] ==1'b1 ? 5'd0 :  
        temp_y[29][9] ==1'b1 ? 5'd31 : 
        temp_y[29][3]==1'b1 ? temp_y[29][8:4]+1'b1 : temp_y[29][8:4];
assign temp_y[30] = 
$signed({3'b0,x140}<<<3'd2)+$signed(-{2'b0,x132}<<<3'd1)+$signed({1'b0,x324})+$signed(-{2'b0,x12}<<<3'd1)+$signed(-{1'b0,x204})+$signed(-{2'b0,x205}<<<3'd1)+$signed(-{2'b0,x69}<<<3'd1)+$signed(-{2'b0,x325}<<<3'd1)+$signed(sharing92)+$signed(-sharing93)-$signed(11'd24);
assign y30=temp_y[30][11] ==1'b1 ? 5'd0 :  
        temp_y[30][9] ==1'b1 ? 5'd31 : 
        temp_y[30][3]==1'b1 ? temp_y[30][8:4]+1'b1 : temp_y[30][8:4];
assign temp_y[31] = 
$signed({2'b0,x268}<<<3'd1)+$signed(-{1'b0,x4})+$signed({1'b0,x204})+$signed({3'b0,x269}<<<3'd2)+$signed(-{1'b0,x324})+$signed(-{1'b0,x197})+$signed(-{1'b0,x5})+$signed(-{1'b0,x76})+$signed(-{1'b0,x196})+$signed(-{1'b0,x333})+$signed(-sharing19)-$signed(11'd32);
assign y31=temp_y[31][11] ==1'b1 ? 5'd0 :  
        temp_y[31][9] ==1'b1 ? 5'd31 : 
        temp_y[31][3]==1'b1 ? temp_y[31][8:4]+1'b1 : temp_y[31][8:4];
assign temp_y[32] = 
$signed(-{1'b0,x68})+$signed(-{1'b0,x5})+$signed({3'b0,x325}<<<3'd2)+$signed(-{2'b0,x269}<<<3'd1)+$signed({3'b0,x333}<<<3'd2)+$signed(-{2'b0,x261}<<<3'd1)+$signed(-{1'b0,x13})+$signed(sharing63)-$signed(11'd0);
assign y32=temp_y[32][11] ==1'b1 ? 5'd0 :  
        temp_y[32][9] ==1'b1 ? 5'd31 : 
        temp_y[32][3]==1'b1 ? temp_y[32][8:4]+1'b1 : temp_y[32][8:4];
assign temp_y[33] = 
$signed(-{1'b0,x197})+$signed(-{2'b0,x260}<<<3'd1)+$signed(-{1'b0,x132})+$signed({1'b0,x196})+$signed({3'b0,x77}<<<3'd2)+$signed({2'b0,x325}<<<3'd1)+$signed({1'b0,x261})+$signed(-{3'b0,x333}<<<3'd2)+$signed(-{1'b0,x332})+$signed(sharing79)-$signed(11'd0);
assign y33=temp_y[33][11] ==1'b1 ? 5'd0 :  
        temp_y[33][9] ==1'b1 ? 5'd31 : 
        temp_y[33][3]==1'b1 ? temp_y[33][8:4]+1'b1 : temp_y[33][8:4];
assign temp_y[34] = 
$signed(-{3'b0,x12}<<<3'd2)+$signed(-{2'b0,x196}<<<3'd1)+$signed({1'b0,x332})+$signed(-{1'b0,x140})+$signed(-{1'b0,x268})+$signed({2'b0,x197}<<<3'd1)+$signed(-{2'b0,x13}<<<3'd1)+$signed(-{2'b0,x141}<<<3'd1)+$signed(-{2'b0,x4}<<<3'd1)+$signed({1'b0,x68})+$signed(sharing31)+$signed(11'd40);
assign y34=temp_y[34][11] ==1'b1 ? 5'd0 :  
        temp_y[34][9] ==1'b1 ? 5'd31 : 
        temp_y[34][3]==1'b1 ? temp_y[34][8:4]+1'b1 : temp_y[34][8:4];
assign temp_y[35] = 
$signed(-{1'b0,x197})+$signed(-{2'b0,x12}<<<3'd1)+$signed({1'b0,x196})+$signed({4'b0,x13}<<<3'd3)+$signed(-{2'b0,x4}<<<3'd1)+$signed(-{2'b0,x205}<<<3'd1)+$signed(-{1'b0,x333})+$signed({1'b0,x68})+$signed(-sharing31)-$signed(11'd8);
assign y35=temp_y[35][11] ==1'b1 ? 5'd0 :  
        temp_y[35][9] ==1'b1 ? 5'd31 : 
        temp_y[35][3]==1'b1 ? temp_y[35][8:4]+1'b1 : temp_y[35][8:4];
assign temp_y[36] = 
$signed({1'b0,x141})+$signed(-{1'b0,x76})+$signed({3'b0,x324}<<<3'd2)+$signed(-{2'b0,x4}<<<3'd1)+$signed(-{1'b0,x12})+$signed({3'b0,x332}<<<3'd2)+$signed(-{1'b0,x268})+$signed({2'b0,x13}<<<3'd1)+$signed(-{1'b0,x69})+$signed({2'b0,x133}<<<3'd1)+$signed(-{1'b0,x140})+$signed(-{2'b0,x204}<<<3'd1)+$signed(-{1'b0,x261})+$signed(-{2'b0,x269}<<<3'd1)+$signed(-{1'b0,x77})+$signed(-{1'b0,x196})+$signed(sharing19)-$signed(11'd16);
assign y36=temp_y[36][11] ==1'b1 ? 5'd0 :  
        temp_y[36][9] ==1'b1 ? 5'd31 : 
        temp_y[36][3]==1'b1 ? temp_y[36][8:4]+1'b1 : temp_y[36][8:4];
assign temp_y[37] = 
$signed(-{1'b0,x197})+$signed(-{1'b0,x323})+$signed(-{4'b0,x268}<<<3'd3)+$signed(-{3'b0,x196}<<<3'd2)+$signed(-{3'b0,x260}<<<3'd2)+$signed(-{1'b0,x331})+$signed(-{4'b0,x261}<<<3'd3)+$signed(-{1'b0,x204})+$signed(-{4'b0,x205}<<<3'd3)+$signed({1'b0,x13})+$signed(-{1'b0,x332})+$signed(-{1'b0,x77})+$signed(-sharing79)+$signed(11'd24);
assign y37=temp_y[37][11] ==1'b1 ? 5'd0 :  
        temp_y[37][9] ==1'b1 ? 5'd31 : 
        temp_y[37][3]==1'b1 ? temp_y[37][8:4]+1'b1 : temp_y[37][8:4];
assign temp_y[38] = 
$signed({1'b0,x68})+$signed({3'b0,x204}<<<3'd2)+$signed({2'b0,x132}<<<3'd1)+$signed({2'b0,x324}<<<3'd1)+$signed(-{2'b0,x268}<<<3'd1)+$signed({1'b0,x332})+$signed(-{1'b0,x12})+$signed(-{3'b0,x133}<<<3'd2)+$signed(-{3'b0,x141}<<<3'd2)+$signed(-{1'b0,x261})+$signed(-{2'b0,x69}<<<3'd1)+$signed({1'b0,x13})+$signed(-{1'b0,x325})+$signed(sharing63)+$signed(11'd16);
assign y38=temp_y[38][11] ==1'b1 ? 5'd0 :  
        temp_y[38][9] ==1'b1 ? 5'd31 : 
        temp_y[38][3]==1'b1 ? temp_y[38][8:4]+1'b1 : temp_y[38][8:4];
assign temp_y[39] = 
$signed({2'b0,x270}<<<3'd1)+$signed(-{1'b0,x79})+$signed(-{3'b0,x335}<<<3'd2)+$signed({1'b0,x142})+$signed(-{3'b0,x334}<<<3'd2)+$signed(-{2'b0,x326}<<<3'd1)+$signed(-{1'b0,x78})+$signed({1'b0,x271})+$signed({2'b0,x263}<<<3'd1)+$signed(-{1'b0,x135})+$signed(sharing48)+$signed(11'd32);
assign y39=temp_y[39][11] ==1'b1 ? 5'd0 :  
        temp_y[39][9] ==1'b1 ? 5'd31 : 
        temp_y[39][3]==1'b1 ? temp_y[39][8:4]+1'b1 : temp_y[39][8:4];
assign temp_y[40] = 
$signed({1'b0,x6})+$signed({2'b0,x78}<<<3'd1)+$signed(-{1'b0,x7})+$signed({1'b0,x70})+$signed(-{1'b0,x142})+$signed({2'b0,x334}<<<3'd1)+$signed(-{1'b0,x270})+$signed({2'b0,x206}<<<3'd1)+$signed({3'b0,x335}<<<3'd2)+$signed(-{2'b0,x207}<<<3'd1)+$signed(-{1'b0,x263})+$signed(sharing48)-$signed(11'd0);
assign y40=temp_y[40][11] ==1'b1 ? 5'd0 :  
        temp_y[40][9] ==1'b1 ? 5'd31 : 
        temp_y[40][3]==1'b1 ? temp_y[40][8:4]+1'b1 : temp_y[40][8:4];
assign temp_y[41] = 
$signed({1'b0,x198})+$signed(-{3'b0,x334}<<<3'd2)+$signed(-{2'b0,x70}<<<3'd1)+$signed(-{2'b0,x78}<<<3'd1)+$signed(-{4'b0,x263}<<<3'd3)+$signed(-{1'b0,x143})+$signed(-{3'b0,x270}<<<3'd2)+$signed(-{2'b0,x326}<<<3'd1)+$signed({1'b0,x134})+$signed({2'b0,x206}<<<3'd1)+$signed(-{3'b0,x271}<<<3'd2)+$signed(-{3'b0,x262}<<<3'd2)+$signed(-{1'b0,x207})+$signed(11'd40);
assign y41=temp_y[41][11] ==1'b1 ? 5'd0 :  
        temp_y[41][9] ==1'b1 ? 5'd31 : 
        temp_y[41][3]==1'b1 ? temp_y[41][8:4]+1'b1 : temp_y[41][8:4];
assign temp_y[42] = 
$signed(-{1'b0,x198})+$signed({1'b0,x327})+$signed({1'b0,x262})+$signed({1'b0,x14})+$signed(-{1'b0,x78})+$signed({1'b0,x142})+$signed({2'b0,x326}<<<3'd1)+$signed(-{1'b0,x70})+$signed(-{2'b0,x79}<<<3'd1)+$signed({1'b0,x271})+$signed(sharing68)+$signed(sharing69)-$signed(11'd16);
assign y42=temp_y[42][11] ==1'b1 ? 5'd0 :  
        temp_y[42][9] ==1'b1 ? 5'd31 : 
        temp_y[42][3]==1'b1 ? temp_y[42][8:4]+1'b1 : temp_y[42][8:4];
assign temp_y[43] = 
$signed(-{2'b0,x14}<<<3'd1)+$signed({1'b0,x326})+$signed({3'b0,x142}<<<3'd2)+$signed(-{2'b0,x134}<<<3'd1)+$signed(-{1'b0,x206})+$signed(-{2'b0,x327}<<<3'd1)+$signed(-{2'b0,x207}<<<3'd1)+$signed(-{2'b0,x71}<<<3'd1)+$signed(sharing68)+$signed(-sharing69)-$signed(11'd24);
assign y43=temp_y[43][11] ==1'b1 ? 5'd0 :  
        temp_y[43][9] ==1'b1 ? 5'd31 : 
        temp_y[43][3]==1'b1 ? temp_y[43][8:4]+1'b1 : temp_y[43][8:4];
assign temp_y[44] = 
$signed(-{1'b0,x198})+$signed({1'b0,x206})+$signed(-{1'b0,x335})+$signed(-{1'b0,x6})+$signed(-{1'b0,x78})+$signed({2'b0,x270}<<<3'd1)+$signed(-{1'b0,x326})+$signed(-{1'b0,x7})+$signed({3'b0,x271}<<<3'd2)+$signed(-{1'b0,x199})+$signed(-sharing25)-$signed(11'd32);
assign y44=temp_y[44][11] ==1'b1 ? 5'd0 :  
        temp_y[44][9] ==1'b1 ? 5'd31 : 
        temp_y[44][3]==1'b1 ? temp_y[44][8:4]+1'b1 : temp_y[44][8:4];
assign temp_y[45] = 
$signed(-{1'b0,x15})+$signed(-{2'b0,x263}<<<3'd1)+$signed({3'b0,x327}<<<3'd2)+$signed(-{1'b0,x70})+$signed({3'b0,x335}<<<3'd2)+$signed(-{2'b0,x271}<<<3'd1)+$signed(-{1'b0,x7})+$signed(sharing56)-$signed(11'd0);
assign y45=temp_y[45][11] ==1'b1 ? 5'd0 :  
        temp_y[45][9] ==1'b1 ? 5'd31 : 
        temp_y[45][3]==1'b1 ? temp_y[45][8:4]+1'b1 : temp_y[45][8:4];
assign temp_y[46] = 
$signed(-{3'b0,x335}<<<3'd2)+$signed(-{1'b0,x334})+$signed(-{1'b0,x199})+$signed(-{1'b0,x134})+$signed(-{2'b0,x262}<<<3'd1)+$signed({1'b0,x198})+$signed({3'b0,x79}<<<3'd2)+$signed({2'b0,x327}<<<3'd1)+$signed({1'b0,x263})+$signed(-sharing96)-$signed(11'd0);
assign y46=temp_y[46][11] ==1'b1 ? 5'd0 :  
        temp_y[46][9] ==1'b1 ? 5'd31 : 
        temp_y[46][3]==1'b1 ? temp_y[46][8:4]+1'b1 : temp_y[46][8:4];
assign temp_y[47] = 
$signed(-{2'b0,x6}<<<3'd1)+$signed(-{2'b0,x143}<<<3'd1)+$signed(-{1'b0,x270})+$signed({2'b0,x199}<<<3'd1)+$signed({1'b0,x70})+$signed({1'b0,x334})+$signed(-{3'b0,x14}<<<3'd2)+$signed(-{2'b0,x198}<<<3'd1)+$signed(-{1'b0,x142})+$signed(-{2'b0,x15}<<<3'd1)+$signed(-sharing6)+$signed(11'd40);
assign y47=temp_y[47][11] ==1'b1 ? 5'd0 :  
        temp_y[47][9] ==1'b1 ? 5'd31 : 
        temp_y[47][3]==1'b1 ? temp_y[47][8:4]+1'b1 : temp_y[47][8:4];
assign temp_y[48] = 
$signed(-{2'b0,x6}<<<3'd1)+$signed({1'b0,x70})+$signed(-{1'b0,x199})+$signed(-{2'b0,x14}<<<3'd1)+$signed({1'b0,x198})+$signed({4'b0,x15}<<<3'd3)+$signed(-{2'b0,x207}<<<3'd1)+$signed(-{1'b0,x335})+$signed(sharing6)-$signed(11'd8);
assign y48=temp_y[48][11] ==1'b1 ? 5'd0 :  
        temp_y[48][9] ==1'b1 ? 5'd31 : 
        temp_y[48][3]==1'b1 ? temp_y[48][8:4]+1'b1 : temp_y[48][8:4];
assign temp_y[49] = 
$signed(-{1'b0,x198})+$signed(-{1'b0,x71})+$signed({3'b0,x326}<<<3'd2)+$signed(-{1'b0,x14})+$signed(-{2'b0,x206}<<<3'd1)+$signed({1'b0,x143})+$signed(-{1'b0,x78})+$signed({2'b0,x15}<<<3'd1)+$signed(-{1'b0,x142})+$signed(-{2'b0,x271}<<<3'd1)+$signed({3'b0,x334}<<<3'd2)+$signed(-{2'b0,x6}<<<3'd1)+$signed(-{1'b0,x270})+$signed(-{1'b0,x263})+$signed({2'b0,x135}<<<3'd1)+$signed(-{1'b0,x79})+$signed(sharing25)-$signed(11'd16);
assign y49=temp_y[49][11] ==1'b1 ? 5'd0 :  
        temp_y[49][9] ==1'b1 ? 5'd31 : 
        temp_y[49][3]==1'b1 ? temp_y[49][8:4]+1'b1 : temp_y[49][8:4];
assign temp_y[50] = 
$signed(-{4'b0,x207}<<<3'd3)+$signed(-{1'b0,x334})+$signed({1'b0,x15})+$signed(-{1'b0,x199})+$signed(-{1'b0,x325})+$signed(-{4'b0,x270}<<<3'd3)+$signed(-{3'b0,x198}<<<3'd2)+$signed(-{1'b0,x206})+$signed(-{4'b0,x263}<<<3'd3)+$signed(-{1'b0,x333})+$signed(-{3'b0,x262}<<<3'd2)+$signed(-{1'b0,x79})+$signed(sharing96)+$signed(11'd24);
assign y50=temp_y[50][11] ==1'b1 ? 5'd0 :  
        temp_y[50][9] ==1'b1 ? 5'd31 : 
        temp_y[50][3]==1'b1 ? temp_y[50][8:4]+1'b1 : temp_y[50][8:4];
assign temp_y[51] = 
$signed(-{3'b0,x143}<<<3'd2)+$signed(-{2'b0,x270}<<<3'd1)+$signed({2'b0,x326}<<<3'd1)+$signed({1'b0,x70})+$signed({1'b0,x334})+$signed({1'b0,x15})+$signed({3'b0,x206}<<<3'd2)+$signed({2'b0,x134}<<<3'd1)+$signed(-{1'b0,x14})+$signed(-{1'b0,x263})+$signed(-{3'b0,x135}<<<3'd2)+$signed(-{2'b0,x71}<<<3'd1)+$signed(-{1'b0,x327})+$signed(sharing56)+$signed(11'd16);
assign y51=temp_y[51][11] ==1'b1 ? 5'd0 :  
        temp_y[51][9] ==1'b1 ? 5'd31 : 
        temp_y[51][3]==1'b1 ? temp_y[51][8:4]+1'b1 : temp_y[51][8:4];
assign temp_y[52] = 
$signed(-{3'b0,x344}<<<3'd2)+$signed({2'b0,x280}<<<3'd1)+$signed(-{1'b0,x88})+$signed(-{2'b0,x336}<<<3'd1)+$signed({1'b0,x152})+$signed({2'b0,x273}<<<3'd1)+$signed({1'b0,x281})+$signed(-{1'b0,x145})+$signed(-{1'b0,x89})+$signed(-{3'b0,x345}<<<3'd2)+$signed(sharing39)+$signed(11'd32);
assign y52=temp_y[52][11] ==1'b1 ? 5'd0 :  
        temp_y[52][9] ==1'b1 ? 5'd31 : 
        temp_y[52][3]==1'b1 ? temp_y[52][8:4]+1'b1 : temp_y[52][8:4];
assign temp_y[53] = 
$signed({2'b0,x344}<<<3'd1)+$signed({1'b0,x16})+$signed({1'b0,x80})+$signed({2'b0,x88}<<<3'd1)+$signed({2'b0,x216}<<<3'd1)+$signed(-{1'b0,x280})+$signed(-{1'b0,x17})+$signed(-{2'b0,x217}<<<3'd1)+$signed(-{1'b0,x273})+$signed(-{1'b0,x152})+$signed({3'b0,x345}<<<3'd2)+$signed(sharing39)-$signed(11'd0);
assign y53=temp_y[53][11] ==1'b1 ? 5'd0 :  
        temp_y[53][9] ==1'b1 ? 5'd31 : 
        temp_y[53][3]==1'b1 ? temp_y[53][8:4]+1'b1 : temp_y[53][8:4];
assign temp_y[54] = 
$signed(-{3'b0,x272}<<<3'd2)+$signed({2'b0,x216}<<<3'd1)+$signed({1'b0,x144})+$signed({1'b0,x208})+$signed(-{2'b0,x80}<<<3'd1)+$signed(-{2'b0,x88}<<<3'd1)+$signed(-{4'b0,x273}<<<3'd3)+$signed(-{3'b0,x280}<<<3'd2)+$signed(-{3'b0,x281}<<<3'd2)+$signed(-{1'b0,x217})+$signed(-{1'b0,x153})+$signed(-{3'b0,x344}<<<3'd2)+$signed(-{2'b0,x336}<<<3'd1)+$signed(11'd40);
assign y54=temp_y[54][11] ==1'b1 ? 5'd0 :  
        temp_y[54][9] ==1'b1 ? 5'd31 : 
        temp_y[54][3]==1'b1 ? temp_y[54][8:4]+1'b1 : temp_y[54][8:4];
assign temp_y[55] = 
$signed({2'b0,x336}<<<3'd1)+$signed({1'b0,x152})+$signed(-{1'b0,x88})+$signed({1'b0,x24})+$signed({1'b0,x272})+$signed({1'b0,x281})+$signed({1'b0,x337})+$signed(-{1'b0,x208})+$signed(-{1'b0,x80})+$signed(-{2'b0,x89}<<<3'd1)+$signed(sharing76)+$signed(-sharing77)-$signed(11'd16);
assign y55=temp_y[55][11] ==1'b1 ? 5'd0 :  
        temp_y[55][9] ==1'b1 ? 5'd31 : 
        temp_y[55][3]==1'b1 ? temp_y[55][8:4]+1'b1 : temp_y[55][8:4];
assign temp_y[56] = 
$signed({3'b0,x152}<<<3'd2)+$signed(-{2'b0,x24}<<<3'd1)+$signed(-{1'b0,x216})+$signed({1'b0,x336})+$signed(-{2'b0,x144}<<<3'd1)+$signed(-{2'b0,x217}<<<3'd1)+$signed(-{2'b0,x81}<<<3'd1)+$signed(-{2'b0,x337}<<<3'd1)+$signed(sharing76)+$signed(sharing77)-$signed(11'd24);
assign y56=temp_y[56][11] ==1'b1 ? 5'd0 :  
        temp_y[56][9] ==1'b1 ? 5'd31 : 
        temp_y[56][3]==1'b1 ? temp_y[56][8:4]+1'b1 : temp_y[56][8:4];
assign temp_y[57] = 
$signed({2'b0,x280}<<<3'd1)+$signed(-{1'b0,x16})+$signed({1'b0,x216})+$signed(-{1'b0,x336})+$signed({3'b0,x281}<<<3'd2)+$signed(-{1'b0,x17})+$signed(-{1'b0,x345})+$signed(-{1'b0,x209})+$signed(-{1'b0,x88})+$signed(-{1'b0,x208})+$signed(sharing27)-$signed(11'd32);
assign y57=temp_y[57][11] ==1'b1 ? 5'd0 :  
        temp_y[57][9] ==1'b1 ? 5'd31 : 
        temp_y[57][3]==1'b1 ? temp_y[57][8:4]+1'b1 : temp_y[57][8:4];
assign temp_y[58] = 
$signed(-{1'b0,x80})+$signed({3'b0,x337}<<<3'd2)+$signed(-{2'b0,x281}<<<3'd1)+$signed({3'b0,x345}<<<3'd2)+$signed(-{2'b0,x273}<<<3'd1)+$signed(-{1'b0,x17})+$signed(-{1'b0,x25})+$signed(sharing62)-$signed(11'd0);
assign y58=temp_y[58][11] ==1'b1 ? 5'd0 :  
        temp_y[58][9] ==1'b1 ? 5'd31 : 
        temp_y[58][3]==1'b1 ? temp_y[58][8:4]+1'b1 : temp_y[58][8:4];
assign temp_y[59] = 
$signed(-{2'b0,x272}<<<3'd1)+$signed(-{1'b0,x144})+$signed({1'b0,x208})+$signed({3'b0,x89}<<<3'd2)+$signed({2'b0,x337}<<<3'd1)+$signed({1'b0,x273})+$signed(-{3'b0,x345}<<<3'd2)+$signed(-{1'b0,x209})+$signed(-{1'b0,x344})+$signed(sharing78)-$signed(11'd0);
assign y59=temp_y[59][11] ==1'b1 ? 5'd0 :  
        temp_y[59][9] ==1'b1 ? 5'd31 : 
        temp_y[59][3]==1'b1 ? temp_y[59][8:4]+1'b1 : temp_y[59][8:4];
assign temp_y[60] = 
$signed(-{3'b0,x24}<<<3'd2)+$signed(-{2'b0,x208}<<<3'd1)+$signed(-{1'b0,x152})+$signed({1'b0,x344})+$signed(-{1'b0,x280})+$signed({2'b0,x209}<<<3'd1)+$signed(-{2'b0,x25}<<<3'd1)+$signed(-{2'b0,x153}<<<3'd1)+$signed(-{2'b0,x16}<<<3'd1)+$signed({1'b0,x80})+$signed(sharing20)+$signed(11'd40);
assign y60=temp_y[60][11] ==1'b1 ? 5'd0 :  
        temp_y[60][9] ==1'b1 ? 5'd31 : 
        temp_y[60][3]==1'b1 ? temp_y[60][8:4]+1'b1 : temp_y[60][8:4];
assign temp_y[61] = 
$signed(-{2'b0,x24}<<<3'd1)+$signed({1'b0,x208})+$signed({4'b0,x25}<<<3'd3)+$signed(-{2'b0,x16}<<<3'd1)+$signed(-{2'b0,x217}<<<3'd1)+$signed(-{1'b0,x345})+$signed(-{1'b0,x209})+$signed({1'b0,x80})+$signed(-sharing20)-$signed(11'd8);
assign y61=temp_y[61][11] ==1'b1 ? 5'd0 :  
        temp_y[61][9] ==1'b1 ? 5'd31 : 
        temp_y[61][3]==1'b1 ? temp_y[61][8:4]+1'b1 : temp_y[61][8:4];
assign temp_y[62] = 
$signed({3'b0,x336}<<<3'd2)+$signed(-{2'b0,x16}<<<3'd1)+$signed(-{1'b0,x24})+$signed(-{1'b0,x152})+$signed({3'b0,x344}<<<3'd2)+$signed({2'b0,x25}<<<3'd1)+$signed({1'b0,x153})+$signed({2'b0,x145}<<<3'd1)+$signed(-{2'b0,x216}<<<3'd1)+$signed(-{2'b0,x281}<<<3'd1)+$signed(-{1'b0,x81})+$signed(-{1'b0,x89})+$signed(-{1'b0,x273})+$signed(-{1'b0,x208})+$signed(-{1'b0,x280})+$signed(-{1'b0,x88})+$signed(-sharing27)-$signed(11'd16);
assign y62=temp_y[62][11] ==1'b1 ? 5'd0 :  
        temp_y[62][9] ==1'b1 ? 5'd31 : 
        temp_y[62][3]==1'b1 ? temp_y[62][8:4]+1'b1 : temp_y[62][8:4];
assign temp_y[63] = 
$signed(-{4'b0,x280}<<<3'd3)+$signed(-{3'b0,x272}<<<3'd2)+$signed(-{3'b0,x208}<<<3'd2)+$signed(-{1'b0,x216})+$signed(-{4'b0,x273}<<<3'd3)+$signed(-{4'b0,x217}<<<3'd3)+$signed(-{1'b0,x335})+$signed({1'b0,x25})+$signed(-{1'b0,x89})+$signed(-{1'b0,x209})+$signed(-{1'b0,x344})+$signed(-{1'b0,x343})+$signed(-sharing78)+$signed(11'd24);
assign y63=temp_y[63][11] ==1'b1 ? 5'd0 :  
        temp_y[63][9] ==1'b1 ? 5'd31 : 
        temp_y[63][3]==1'b1 ? temp_y[63][8:4]+1'b1 : temp_y[63][8:4];
assign temp_y[64] = 
$signed({3'b0,x216}<<<3'd2)+$signed({2'b0,x144}<<<3'd1)+$signed({1'b0,x344})+$signed({2'b0,x336}<<<3'd1)+$signed(-{2'b0,x280}<<<3'd1)+$signed(-{1'b0,x24})+$signed(-{3'b0,x153}<<<3'd2)+$signed(-{3'b0,x145}<<<3'd2)+$signed(-{2'b0,x81}<<<3'd1)+$signed(-{1'b0,x273})+$signed(-{1'b0,x337})+$signed({1'b0,x25})+$signed({1'b0,x80})+$signed(sharing62)+$signed(11'd16);
assign y64=temp_y[64][11] ==1'b1 ? 5'd0 :  
        temp_y[64][9] ==1'b1 ? 5'd31 : 
        temp_y[64][3]==1'b1 ? temp_y[64][8:4]+1'b1 : temp_y[64][8:4];
assign temp_y[65] = 
$signed(-{3'b0,x346}<<<3'd2)+$signed({2'b0,x282}<<<3'd1)+$signed(-{1'b0,x90})+$signed(-{2'b0,x338}<<<3'd1)+$signed({1'b0,x154})+$signed({2'b0,x275}<<<3'd1)+$signed({1'b0,x283})+$signed(-{1'b0,x147})+$signed(-{1'b0,x91})+$signed(-{3'b0,x347}<<<3'd2)+$signed(sharing46)+$signed(11'd32);
assign y65=temp_y[65][11] ==1'b1 ? 5'd0 :  
        temp_y[65][9] ==1'b1 ? 5'd31 : 
        temp_y[65][3]==1'b1 ? temp_y[65][8:4]+1'b1 : temp_y[65][8:4];
assign temp_y[66] = 
$signed({2'b0,x218}<<<3'd1)+$signed({1'b0,x82})+$signed({1'b0,x18})+$signed({2'b0,x346}<<<3'd1)+$signed({2'b0,x90}<<<3'd1)+$signed(-{1'b0,x282})+$signed(-{1'b0,x19})+$signed(-{2'b0,x219}<<<3'd1)+$signed(-{1'b0,x275})+$signed(-{1'b0,x154})+$signed({3'b0,x347}<<<3'd2)+$signed(sharing46)-$signed(11'd0);
assign y66=temp_y[66][11] ==1'b1 ? 5'd0 :  
        temp_y[66][9] ==1'b1 ? 5'd31 : 
        temp_y[66][3]==1'b1 ? temp_y[66][8:4]+1'b1 : temp_y[66][8:4];
assign temp_y[67] = 
$signed(-{3'b0,x274}<<<3'd2)+$signed({2'b0,x218}<<<3'd1)+$signed({1'b0,x146})+$signed({1'b0,x210})+$signed(-{2'b0,x82}<<<3'd1)+$signed(-{2'b0,x90}<<<3'd1)+$signed(-{4'b0,x275}<<<3'd3)+$signed(-{3'b0,x282}<<<3'd2)+$signed(-{3'b0,x283}<<<3'd2)+$signed(-{1'b0,x219})+$signed(-{1'b0,x155})+$signed(-{3'b0,x346}<<<3'd2)+$signed(-{2'b0,x338}<<<3'd1)+$signed(11'd40);
assign y67=temp_y[67][11] ==1'b1 ? 5'd0 :  
        temp_y[67][9] ==1'b1 ? 5'd31 : 
        temp_y[67][3]==1'b1 ? temp_y[67][8:4]+1'b1 : temp_y[67][8:4];
assign temp_y[68] = 
$signed({2'b0,x338}<<<3'd1)+$signed({1'b0,x154})+$signed({1'b0,x26})+$signed({1'b0,x274})+$signed(-{1'b0,x90})+$signed({1'b0,x339})+$signed({1'b0,x283})+$signed(-{1'b0,x210})+$signed(-{1'b0,x82})+$signed(-{2'b0,x91}<<<3'd1)+$signed(sharing101)+$signed(sharing102)-$signed(11'd16);
assign y68=temp_y[68][11] ==1'b1 ? 5'd0 :  
        temp_y[68][9] ==1'b1 ? 5'd31 : 
        temp_y[68][3]==1'b1 ? temp_y[68][8:4]+1'b1 : temp_y[68][8:4];
assign temp_y[69] = 
$signed({3'b0,x154}<<<3'd2)+$signed(-{2'b0,x26}<<<3'd1)+$signed(-{1'b0,x218})+$signed({1'b0,x338})+$signed(-{2'b0,x146}<<<3'd1)+$signed(-{2'b0,x219}<<<3'd1)+$signed(-{2'b0,x83}<<<3'd1)+$signed(-{2'b0,x339}<<<3'd1)+$signed(sharing101)+$signed(-sharing102)-$signed(11'd24);
assign y69=temp_y[69][11] ==1'b1 ? 5'd0 :  
        temp_y[69][9] ==1'b1 ? 5'd31 : 
        temp_y[69][3]==1'b1 ? temp_y[69][8:4]+1'b1 : temp_y[69][8:4];
assign temp_y[70] = 
$signed({2'b0,x282}<<<3'd1)+$signed(-{1'b0,x18})+$signed({1'b0,x218})+$signed(-{1'b0,x338})+$signed({3'b0,x283}<<<3'd2)+$signed(-{1'b0,x211})+$signed(-{1'b0,x19})+$signed(-{1'b0,x347})+$signed(-{1'b0,x90})+$signed(-{1'b0,x210})+$signed(-sharing24)-$signed(11'd32);
assign y70=temp_y[70][11] ==1'b1 ? 5'd0 :  
        temp_y[70][9] ==1'b1 ? 5'd31 : 
        temp_y[70][3]==1'b1 ? temp_y[70][8:4]+1'b1 : temp_y[70][8:4];
assign temp_y[71] = 
$signed(-{1'b0,x82})+$signed({3'b0,x347}<<<3'd2)+$signed(-{2'b0,x275}<<<3'd1)+$signed({3'b0,x339}<<<3'd2)+$signed(-{2'b0,x283}<<<3'd1)+$signed(-{1'b0,x19})+$signed(-{1'b0,x27})+$signed(sharing55)-$signed(11'd0);
assign y71=temp_y[71][11] ==1'b1 ? 5'd0 :  
        temp_y[71][9] ==1'b1 ? 5'd31 : 
        temp_y[71][3]==1'b1 ? temp_y[71][8:4]+1'b1 : temp_y[71][8:4];
assign temp_y[72] = 
$signed(-{2'b0,x274}<<<3'd1)+$signed({1'b0,x210})+$signed(-{1'b0,x146})+$signed({3'b0,x91}<<<3'd2)+$signed(-{3'b0,x347}<<<3'd2)+$signed({2'b0,x339}<<<3'd1)+$signed({1'b0,x275})+$signed(-{1'b0,x211})+$signed(-{1'b0,x346})+$signed(sharing100)-$signed(11'd0);
assign y72=temp_y[72][11] ==1'b1 ? 5'd0 :  
        temp_y[72][9] ==1'b1 ? 5'd31 : 
        temp_y[72][3]==1'b1 ? temp_y[72][8:4]+1'b1 : temp_y[72][8:4];
assign temp_y[73] = 
$signed(-{3'b0,x26}<<<3'd2)+$signed(-{2'b0,x210}<<<3'd1)+$signed(-{1'b0,x154})+$signed({1'b0,x346})+$signed(-{1'b0,x282})+$signed({2'b0,x211}<<<3'd1)+$signed(-{2'b0,x27}<<<3'd1)+$signed(-{2'b0,x155}<<<3'd1)+$signed(-{2'b0,x18}<<<3'd1)+$signed({1'b0,x82})+$signed(sharing5)+$signed(11'd40);
assign y73=temp_y[73][11] ==1'b1 ? 5'd0 :  
        temp_y[73][9] ==1'b1 ? 5'd31 : 
        temp_y[73][3]==1'b1 ? temp_y[73][8:4]+1'b1 : temp_y[73][8:4];
assign temp_y[74] = 
$signed(-{2'b0,x26}<<<3'd1)+$signed({1'b0,x210})+$signed({4'b0,x27}<<<3'd3)+$signed(-{2'b0,x18}<<<3'd1)+$signed(-{2'b0,x219}<<<3'd1)+$signed(-{1'b0,x211})+$signed(-{1'b0,x347})+$signed({1'b0,x82})+$signed(-sharing5)-$signed(11'd8);
assign y74=temp_y[74][11] ==1'b1 ? 5'd0 :  
        temp_y[74][9] ==1'b1 ? 5'd31 : 
        temp_y[74][3]==1'b1 ? temp_y[74][8:4]+1'b1 : temp_y[74][8:4];
assign temp_y[75] = 
$signed(-{1'b0,x90})+$signed({3'b0,x338}<<<3'd2)+$signed(-{2'b0,x18}<<<3'd1)+$signed(-{1'b0,x26})+$signed(-{1'b0,x154})+$signed({3'b0,x346}<<<3'd2)+$signed({2'b0,x27}<<<3'd1)+$signed({1'b0,x155})+$signed({2'b0,x147}<<<3'd1)+$signed(-{2'b0,x218}<<<3'd1)+$signed(-{2'b0,x283}<<<3'd1)+$signed(-{1'b0,x83})+$signed(-{1'b0,x91})+$signed(-{1'b0,x275})+$signed(-{1'b0,x210})+$signed(-{1'b0,x282})+$signed(sharing24)-$signed(11'd16);
assign y75=temp_y[75][11] ==1'b1 ? 5'd0 :  
        temp_y[75][9] ==1'b1 ? 5'd31 : 
        temp_y[75][3]==1'b1 ? temp_y[75][8:4]+1'b1 : temp_y[75][8:4];
assign temp_y[76] = 
$signed(-{1'b0,x337})+$signed(-{4'b0,x282}<<<3'd3)+$signed(-{3'b0,x210}<<<3'd2)+$signed(-{3'b0,x274}<<<3'd2)+$signed(-{1'b0,x345})+$signed(-{4'b0,x275}<<<3'd3)+$signed(-{1'b0,x218})+$signed(-{4'b0,x219}<<<3'd3)+$signed({1'b0,x27})+$signed(-{1'b0,x91})+$signed(-{1'b0,x211})+$signed(-{1'b0,x346})+$signed(-sharing100)+$signed(11'd24);
assign y76=temp_y[76][11] ==1'b1 ? 5'd0 :  
        temp_y[76][9] ==1'b1 ? 5'd31 : 
        temp_y[76][3]==1'b1 ? temp_y[76][8:4]+1'b1 : temp_y[76][8:4];
assign temp_y[77] = 
$signed({1'b0,x82})+$signed({3'b0,x218}<<<3'd2)+$signed({2'b0,x146}<<<3'd1)+$signed({1'b0,x346})+$signed({2'b0,x338}<<<3'd1)+$signed(-{3'b0,x147}<<<3'd2)+$signed(-{2'b0,x282}<<<3'd1)+$signed(-{1'b0,x339})+$signed(-{1'b0,x26})+$signed(-{3'b0,x155}<<<3'd2)+$signed(-{2'b0,x83}<<<3'd1)+$signed(-{1'b0,x275})+$signed({1'b0,x27})+$signed(sharing55)+$signed(11'd16);
assign y77=temp_y[77][11] ==1'b1 ? 5'd0 :  
        temp_y[77][9] ==1'b1 ? 5'd31 : 
        temp_y[77][3]==1'b1 ? temp_y[77][8:4]+1'b1 : temp_y[77][8:4];
assign temp_y[78] = 
$signed(-{3'b0,x348}<<<3'd2)+$signed({2'b0,x284}<<<3'd1)+$signed(-{1'b0,x92})+$signed(-{2'b0,x340}<<<3'd1)+$signed({1'b0,x285})+$signed({2'b0,x277}<<<3'd1)+$signed(-{1'b0,x149})+$signed({1'b0,x156})+$signed(-{3'b0,x349}<<<3'd2)+$signed(-{1'b0,x93})+$signed(sharing38)+$signed(11'd32);
assign y78=temp_y[78][11] ==1'b1 ? 5'd0 :  
        temp_y[78][9] ==1'b1 ? 5'd31 : 
        temp_y[78][3]==1'b1 ? temp_y[78][8:4]+1'b1 : temp_y[78][8:4];
assign temp_y[79] = 
$signed({2'b0,x348}<<<3'd1)+$signed({1'b0,x20})+$signed({1'b0,x84})+$signed({2'b0,x92}<<<3'd1)+$signed({2'b0,x220}<<<3'd1)+$signed(-{1'b0,x284})+$signed(-{1'b0,x21})+$signed(-{2'b0,x221}<<<3'd1)+$signed(-{1'b0,x277})+$signed(-{1'b0,x156})+$signed({3'b0,x349}<<<3'd2)+$signed(sharing38)-$signed(11'd0);
assign y79=temp_y[79][11] ==1'b1 ? 5'd0 :  
        temp_y[79][9] ==1'b1 ? 5'd31 : 
        temp_y[79][3]==1'b1 ? temp_y[79][8:4]+1'b1 : temp_y[79][8:4];
assign temp_y[80] = 
$signed(-{2'b0,x340}<<<3'd1)+$signed(-{1'b0,x157})+$signed(-{3'b0,x276}<<<3'd2)+$signed(-{3'b0,x348}<<<3'd2)+$signed({2'b0,x220}<<<3'd1)+$signed({1'b0,x212})+$signed({1'b0,x148})+$signed(-{2'b0,x84}<<<3'd1)+$signed(-{1'b0,x221})+$signed(-{2'b0,x92}<<<3'd1)+$signed(-{4'b0,x277}<<<3'd3)+$signed(-{3'b0,x284}<<<3'd2)+$signed(-{3'b0,x285}<<<3'd2)+$signed(11'd40);
assign y80=temp_y[80][11] ==1'b1 ? 5'd0 :  
        temp_y[80][9] ==1'b1 ? 5'd31 : 
        temp_y[80][3]==1'b1 ? temp_y[80][8:4]+1'b1 : temp_y[80][8:4];
assign temp_y[81] = 
$signed({2'b0,x340}<<<3'd1)+$signed({1'b0,x156})+$signed(-{1'b0,x92})+$signed({1'b0,x28})+$signed({1'b0,x276})+$signed({1'b0,x285})+$signed(-{1'b0,x212})+$signed(-{1'b0,x84})+$signed(-{2'b0,x93}<<<3'd1)+$signed({1'b0,x341})+$signed(sharing74)+$signed(sharing75)-$signed(11'd16);
assign y81=temp_y[81][11] ==1'b1 ? 5'd0 :  
        temp_y[81][9] ==1'b1 ? 5'd31 : 
        temp_y[81][3]==1'b1 ? temp_y[81][8:4]+1'b1 : temp_y[81][8:4];
assign temp_y[82] = 
$signed({3'b0,x156}<<<3'd2)+$signed(-{2'b0,x28}<<<3'd1)+$signed(-{1'b0,x220})+$signed({1'b0,x340})+$signed(-{2'b0,x148}<<<3'd1)+$signed(-{2'b0,x221}<<<3'd1)+$signed(-{2'b0,x85}<<<3'd1)+$signed(-{2'b0,x341}<<<3'd1)+$signed(sharing74)+$signed(-sharing75)-$signed(11'd24);
assign y82=temp_y[82][11] ==1'b1 ? 5'd0 :  
        temp_y[82][9] ==1'b1 ? 5'd31 : 
        temp_y[82][3]==1'b1 ? temp_y[82][8:4]+1'b1 : temp_y[82][8:4];
assign temp_y[83] = 
$signed({2'b0,x284}<<<3'd1)+$signed(-{1'b0,x20})+$signed({1'b0,x220})+$signed(-{1'b0,x340})+$signed({3'b0,x285}<<<3'd2)+$signed(-{1'b0,x213})+$signed(-{1'b0,x21})+$signed(-{1'b0,x92})+$signed(-{1'b0,x212})+$signed(-{1'b0,x349})+$signed(-sharing14)-$signed(11'd32);
assign y83=temp_y[83][11] ==1'b1 ? 5'd0 :  
        temp_y[83][9] ==1'b1 ? 5'd31 : 
        temp_y[83][3]==1'b1 ? temp_y[83][8:4]+1'b1 : temp_y[83][8:4];
assign temp_y[84] = 
$signed(-{1'b0,x84})+$signed(-{1'b0,x29})+$signed({3'b0,x341}<<<3'd2)+$signed(-{2'b0,x285}<<<3'd1)+$signed({3'b0,x349}<<<3'd2)+$signed(-{2'b0,x277}<<<3'd1)+$signed(-{1'b0,x21})+$signed(sharing61)-$signed(11'd0);
assign y84=temp_y[84][11] ==1'b1 ? 5'd0 :  
        temp_y[84][9] ==1'b1 ? 5'd31 : 
        temp_y[84][3]==1'b1 ? temp_y[84][8:4]+1'b1 : temp_y[84][8:4];
assign temp_y[85] = 
$signed(-{1'b0,x213})+$signed(-{2'b0,x276}<<<3'd1)+$signed(-{1'b0,x148})+$signed({1'b0,x212})+$signed({3'b0,x93}<<<3'd2)+$signed({2'b0,x341}<<<3'd1)+$signed({1'b0,x277})+$signed(-{3'b0,x349}<<<3'd2)+$signed(-{1'b0,x348})+$signed(-sharing86)-$signed(11'd0);
assign y85=temp_y[85][11] ==1'b1 ? 5'd0 :  
        temp_y[85][9] ==1'b1 ? 5'd31 : 
        temp_y[85][3]==1'b1 ? temp_y[85][8:4]+1'b1 : temp_y[85][8:4];
assign temp_y[86] = 
$signed(-{3'b0,x28}<<<3'd2)+$signed(-{2'b0,x212}<<<3'd1)+$signed(-{1'b0,x156})+$signed({1'b0,x348})+$signed(-{1'b0,x284})+$signed({2'b0,x213}<<<3'd1)+$signed(-{2'b0,x29}<<<3'd1)+$signed(-{2'b0,x157}<<<3'd1)+$signed(-{2'b0,x20}<<<3'd1)+$signed({1'b0,x84})+$signed(sharing17)+$signed(11'd40);
assign y86=temp_y[86][11] ==1'b1 ? 5'd0 :  
        temp_y[86][9] ==1'b1 ? 5'd31 : 
        temp_y[86][3]==1'b1 ? temp_y[86][8:4]+1'b1 : temp_y[86][8:4];
assign temp_y[87] = 
$signed(-{1'b0,x213})+$signed(-{2'b0,x28}<<<3'd1)+$signed({1'b0,x212})+$signed({4'b0,x29}<<<3'd3)+$signed(-{2'b0,x20}<<<3'd1)+$signed(-{2'b0,x221}<<<3'd1)+$signed(-{1'b0,x349})+$signed({1'b0,x84})+$signed(-sharing17)-$signed(11'd8);
assign y87=temp_y[87][11] ==1'b1 ? 5'd0 :  
        temp_y[87][9] ==1'b1 ? 5'd31 : 
        temp_y[87][3]==1'b1 ? temp_y[87][8:4]+1'b1 : temp_y[87][8:4];
assign temp_y[88] = 
$signed(-{1'b0,x212})+$signed(-{1'b0,x92})+$signed({3'b0,x340}<<<3'd2)+$signed(-{2'b0,x20}<<<3'd1)+$signed(-{1'b0,x28})+$signed(-{1'b0,x156})+$signed({3'b0,x348}<<<3'd2)+$signed({2'b0,x149}<<<3'd1)+$signed({1'b0,x157})+$signed({2'b0,x29}<<<3'd1)+$signed(-{2'b0,x220}<<<3'd1)+$signed(-{1'b0,x277})+$signed(-{1'b0,x284})+$signed(-{2'b0,x285}<<<3'd1)+$signed(-{1'b0,x85})+$signed(-{1'b0,x93})+$signed(sharing14)-$signed(11'd16);
assign y88=temp_y[88][11] ==1'b1 ? 5'd0 :  
        temp_y[88][9] ==1'b1 ? 5'd31 : 
        temp_y[88][3]==1'b1 ? temp_y[88][8:4]+1'b1 : temp_y[88][8:4];
assign temp_y[89] = 
$signed(-{1'b0,x213})+$signed(-{1'b0,x339})+$signed(-{4'b0,x284}<<<3'd3)+$signed(-{3'b0,x212}<<<3'd2)+$signed(-{3'b0,x276}<<<3'd2)+$signed(-{1'b0,x347})+$signed(-{4'b0,x277}<<<3'd3)+$signed(-{1'b0,x220})+$signed(-{4'b0,x221}<<<3'd3)+$signed({1'b0,x29})+$signed(-{1'b0,x348})+$signed(-{1'b0,x93})+$signed(sharing86)+$signed(11'd24);
assign y89=temp_y[89][11] ==1'b1 ? 5'd0 :  
        temp_y[89][9] ==1'b1 ? 5'd31 : 
        temp_y[89][3]==1'b1 ? temp_y[89][8:4]+1'b1 : temp_y[89][8:4];
assign temp_y[90] = 
$signed({3'b0,x220}<<<3'd2)+$signed({2'b0,x148}<<<3'd1)+$signed({1'b0,x348})+$signed({2'b0,x340}<<<3'd1)+$signed(-{2'b0,x284}<<<3'd1)+$signed(-{1'b0,x28})+$signed(-{3'b0,x157}<<<3'd2)+$signed(-{3'b0,x149}<<<3'd2)+$signed(-{2'b0,x85}<<<3'd1)+$signed(-{1'b0,x277})+$signed({1'b0,x29})+$signed({1'b0,x84})+$signed(-{1'b0,x341})+$signed(sharing61)+$signed(11'd16);
assign y90=temp_y[90][11] ==1'b1 ? 5'd0 :  
        temp_y[90][9] ==1'b1 ? 5'd31 : 
        temp_y[90][3]==1'b1 ? temp_y[90][8:4]+1'b1 : temp_y[90][8:4];
assign temp_y[91] = 
$signed(-{1'b0,x95})+$signed({1'b0,x158})+$signed(-{2'b0,x342}<<<3'd1)+$signed(-{3'b0,x351}<<<3'd2)+$signed(-{3'b0,x350}<<<3'd2)+$signed({2'b0,x286}<<<3'd1)+$signed(-{1'b0,x94})+$signed({1'b0,x287})+$signed({2'b0,x279}<<<3'd1)+$signed(-{1'b0,x151})+$signed(sharing44)+$signed(11'd32);
assign y91=temp_y[91][11] ==1'b1 ? 5'd0 :  
        temp_y[91][9] ==1'b1 ? 5'd31 : 
        temp_y[91][3]==1'b1 ? temp_y[91][8:4]+1'b1 : temp_y[91][8:4];
assign temp_y[92] = 
$signed(-{1'b0,x158})+$signed({1'b0,x22})+$signed({2'b0,x350}<<<3'd1)+$signed({1'b0,x86})+$signed(-{2'b0,x223}<<<3'd1)+$signed(-{1'b0,x279})+$signed({2'b0,x94}<<<3'd1)+$signed(-{1'b0,x286})+$signed({3'b0,x351}<<<3'd2)+$signed({2'b0,x222}<<<3'd1)+$signed(-{1'b0,x23})+$signed(sharing44)-$signed(11'd0);
assign y92=temp_y[92][11] ==1'b1 ? 5'd0 :  
        temp_y[92][9] ==1'b1 ? 5'd31 : 
        temp_y[92][3]==1'b1 ? temp_y[92][8:4]+1'b1 : temp_y[92][8:4];
assign temp_y[93] = 
$signed(-{3'b0,x286}<<<3'd2)+$signed({1'b0,x214})+$signed(-{3'b0,x350}<<<3'd2)+$signed(-{2'b0,x86}<<<3'd1)+$signed(-{2'b0,x94}<<<3'd1)+$signed(-{1'b0,x159})+$signed(-{3'b0,x278}<<<3'd2)+$signed(-{2'b0,x342}<<<3'd1)+$signed({1'b0,x150})+$signed(-{4'b0,x279}<<<3'd3)+$signed(-{3'b0,x287}<<<3'd2)+$signed({2'b0,x222}<<<3'd1)+$signed(-{1'b0,x223})+$signed(11'd40);
assign y93=temp_y[93][11] ==1'b1 ? 5'd0 :  
        temp_y[93][9] ==1'b1 ? 5'd31 : 
        temp_y[93][3]==1'b1 ? temp_y[93][8:4]+1'b1 : temp_y[93][8:4];
assign temp_y[94] = 
$signed(-{1'b0,x214})+$signed({1'b0,x343})+$signed({1'b0,x278})+$signed({1'b0,x30})+$signed(-{1'b0,x86})+$signed(-{1'b0,x94})+$signed({2'b0,x342}<<<3'd1)+$signed({1'b0,x158})+$signed(-{2'b0,x95}<<<3'd1)+$signed({1'b0,x287})+$signed(sharing94)+$signed(sharing95)-$signed(11'd16);
assign y94=temp_y[94][11] ==1'b1 ? 5'd0 :  
        temp_y[94][9] ==1'b1 ? 5'd31 : 
        temp_y[94][3]==1'b1 ? temp_y[94][8:4]+1'b1 : temp_y[94][8:4];
assign temp_y[95] = 
$signed(-{2'b0,x87}<<<3'd1)+$signed(-{2'b0,x343}<<<3'd1)+$signed({1'b0,x342})+$signed(-{2'b0,x150}<<<3'd1)+$signed({3'b0,x158}<<<3'd2)+$signed(-{2'b0,x30}<<<3'd1)+$signed(-{1'b0,x222})+$signed(-{2'b0,x223}<<<3'd1)+$signed(sharing94)+$signed(-sharing95)-$signed(11'd24);
assign y95=temp_y[95][11] ==1'b1 ? 5'd0 :  
        temp_y[95][9] ==1'b1 ? 5'd31 : 
        temp_y[95][3]==1'b1 ? temp_y[95][8:4]+1'b1 : temp_y[95][8:4];
assign temp_y[96] = 
$signed(-{1'b0,x214})+$signed(-{1'b0,x22})+$signed(-{1'b0,x342})+$signed(-{1'b0,x94})+$signed(-{1'b0,x215})+$signed({2'b0,x286}<<<3'd1)+$signed({1'b0,x222})+$signed({3'b0,x287}<<<3'd2)+$signed(-{1'b0,x23})+$signed(-{1'b0,x351})+$signed(sharing11)-$signed(11'd32);
assign y96=temp_y[96][11] ==1'b1 ? 5'd0 :  
        temp_y[96][9] ==1'b1 ? 5'd31 : 
        temp_y[96][3]==1'b1 ? temp_y[96][8:4]+1'b1 : temp_y[96][8:4];
assign temp_y[97] = 
$signed(-{1'b0,x31})+$signed(-{2'b0,x279}<<<3'd1)+$signed(-{1'b0,x86})+$signed({3'b0,x343}<<<3'd2)+$signed({3'b0,x351}<<<3'd2)+$signed(-{2'b0,x287}<<<3'd1)+$signed(-{1'b0,x23})+$signed(sharing57)-$signed(11'd0);
assign y97=temp_y[97][11] ==1'b1 ? 5'd0 :  
        temp_y[97][9] ==1'b1 ? 5'd31 : 
        temp_y[97][3]==1'b1 ? temp_y[97][8:4]+1'b1 : temp_y[97][8:4];
assign temp_y[98] = 
$signed(-{1'b0,x150})+$signed(-{3'b0,x351}<<<3'd2)+$signed(-{1'b0,x350})+$signed(-{1'b0,x215})+$signed(-{2'b0,x278}<<<3'd1)+$signed({1'b0,x214})+$signed({3'b0,x95}<<<3'd2)+$signed({2'b0,x343}<<<3'd1)+$signed({1'b0,x279})+$signed(sharing91)-$signed(11'd0);
assign y98=temp_y[98][11] ==1'b1 ? 5'd0 :  
        temp_y[98][9] ==1'b1 ? 5'd31 : 
        temp_y[98][3]==1'b1 ? temp_y[98][8:4]+1'b1 : temp_y[98][8:4];
assign temp_y[99] = 
$signed(-{2'b0,x22}<<<3'd1)+$signed(-{1'b0,x158})+$signed({2'b0,x215}<<<3'd1)+$signed({1'b0,x86})+$signed({1'b0,x350})+$signed(-{3'b0,x30}<<<3'd2)+$signed(-{2'b0,x31}<<<3'd1)+$signed(-{1'b0,x286})+$signed(-{2'b0,x214}<<<3'd1)+$signed(-{2'b0,x159}<<<3'd1)+$signed(sharing0)+$signed(11'd40);
assign y99=temp_y[99][11] ==1'b1 ? 5'd0 :  
        temp_y[99][9] ==1'b1 ? 5'd31 : 
        temp_y[99][3]==1'b1 ? temp_y[99][8:4]+1'b1 : temp_y[99][8:4];
assign temp_y[100] = 
$signed(-{2'b0,x22}<<<3'd1)+$signed({1'b0,x86})+$signed(-{1'b0,x215})+$signed(-{2'b0,x30}<<<3'd1)+$signed({1'b0,x214})+$signed({4'b0,x31}<<<3'd3)+$signed(-{2'b0,x223}<<<3'd1)+$signed(-{1'b0,x351})+$signed(-sharing0)-$signed(11'd8);
assign y100=temp_y[100][11] ==1'b1 ? 5'd0 :  
        temp_y[100][9] ==1'b1 ? 5'd31 : 
        temp_y[100][3]==1'b1 ? temp_y[100][8:4]+1'b1 : temp_y[100][8:4];
assign temp_y[101] = 
$signed(-{1'b0,x214})+$signed({2'b0,x31}<<<3'd1)+$signed(-{1'b0,x87})+$signed({3'b0,x342}<<<3'd2)+$signed({2'b0,x151}<<<3'd1)+$signed(-{1'b0,x158})+$signed(-{1'b0,x30})+$signed({1'b0,x159})+$signed(-{1'b0,x94})+$signed(-{2'b0,x222}<<<3'd1)+$signed(-{1'b0,x279})+$signed({3'b0,x350}<<<3'd2)+$signed(-{2'b0,x22}<<<3'd1)+$signed(-{1'b0,x286})+$signed(-{2'b0,x287}<<<3'd1)+$signed(-{1'b0,x95})+$signed(-sharing11)-$signed(11'd16);
assign y101=temp_y[101][11] ==1'b1 ? 5'd0 :  
        temp_y[101][9] ==1'b1 ? 5'd31 : 
        temp_y[101][3]==1'b1 ? temp_y[101][8:4]+1'b1 : temp_y[101][8:4];
assign temp_y[102] = 
$signed(-{4'b0,x223}<<<3'd3)+$signed({1'b0,x31})+$signed(-{1'b0,x350})+$signed(-{1'b0,x215})+$signed(-{1'b0,x341})+$signed(-{4'b0,x286}<<<3'd3)+$signed(-{3'b0,x278}<<<3'd2)+$signed(-{1'b0,x222})+$signed(-{4'b0,x279}<<<3'd3)+$signed(-{1'b0,x349})+$signed(-{3'b0,x214}<<<3'd2)+$signed(-{1'b0,x95})+$signed(-sharing91)+$signed(11'd24);
assign y102=temp_y[102][11] ==1'b1 ? 5'd0 :  
        temp_y[102][9] ==1'b1 ? 5'd31 : 
        temp_y[102][3]==1'b1 ? temp_y[102][8:4]+1'b1 : temp_y[102][8:4];
assign temp_y[103] = 
$signed(-{3'b0,x151}<<<3'd2)+$signed(-{2'b0,x286}<<<3'd1)+$signed({1'b0,x86})+$signed({1'b0,x350})+$signed({2'b0,x150}<<<3'd1)+$signed(-{1'b0,x279})+$signed({3'b0,x222}<<<3'd2)+$signed({2'b0,x342}<<<3'd1)+$signed(-{1'b0,x30})+$signed({1'b0,x31})+$signed(-{3'b0,x159}<<<3'd2)+$signed(-{2'b0,x87}<<<3'd1)+$signed(-{1'b0,x343})+$signed(sharing57)+$signed(11'd16);
assign y103=temp_y[103][11] ==1'b1 ? 5'd0 :  
        temp_y[103][9] ==1'b1 ? 5'd31 : 
        temp_y[103][3]==1'b1 ? temp_y[103][8:4]+1'b1 : temp_y[103][8:4];
assign temp_y[104] = 
$signed(-{3'b0,x360}<<<3'd2)+$signed({2'b0,x296}<<<3'd1)+$signed(-{1'b0,x104})+$signed(-{2'b0,x352}<<<3'd1)+$signed({1'b0,x168})+$signed({2'b0,x289}<<<3'd1)+$signed({1'b0,x297})+$signed(-{1'b0,x105})+$signed(-{1'b0,x161})+$signed(-{3'b0,x361}<<<3'd2)+$signed(sharing35)+$signed(11'd32);
assign y104=temp_y[104][11] ==1'b1 ? 5'd0 :  
        temp_y[104][9] ==1'b1 ? 5'd31 : 
        temp_y[104][3]==1'b1 ? temp_y[104][8:4]+1'b1 : temp_y[104][8:4];
assign temp_y[105] = 
$signed({2'b0,x232}<<<3'd1)+$signed({2'b0,x104}<<<3'd1)+$signed({2'b0,x360}<<<3'd1)+$signed({1'b0,x32})+$signed({1'b0,x96})+$signed(-{1'b0,x33})+$signed(-{1'b0,x296})+$signed(-{2'b0,x233}<<<3'd1)+$signed(-{1'b0,x289})+$signed(-{1'b0,x168})+$signed({3'b0,x361}<<<3'd2)+$signed(sharing35)-$signed(11'd0);
assign y105=temp_y[105][11] ==1'b1 ? 5'd0 :  
        temp_y[105][9] ==1'b1 ? 5'd31 : 
        temp_y[105][3]==1'b1 ? temp_y[105][8:4]+1'b1 : temp_y[105][8:4];
assign temp_y[106] = 
$signed(-{3'b0,x288}<<<3'd2)+$signed(-{2'b0,x104}<<<3'd1)+$signed({2'b0,x232}<<<3'd1)+$signed({1'b0,x160})+$signed({1'b0,x224})+$signed(-{2'b0,x96}<<<3'd1)+$signed(-{4'b0,x289}<<<3'd3)+$signed(-{3'b0,x296}<<<3'd2)+$signed(-{3'b0,x297}<<<3'd2)+$signed(-{1'b0,x233})+$signed(-{1'b0,x169})+$signed(-{3'b0,x360}<<<3'd2)+$signed(-{2'b0,x352}<<<3'd1)+$signed(11'd40);
assign y106=temp_y[106][11] ==1'b1 ? 5'd0 :  
        temp_y[106][9] ==1'b1 ? 5'd31 : 
        temp_y[106][3]==1'b1 ? temp_y[106][8:4]+1'b1 : temp_y[106][8:4];
assign temp_y[107] = 
$signed({2'b0,x352}<<<3'd1)+$signed(-{1'b0,x96})+$signed({1'b0,x40})+$signed({1'b0,x288})+$signed({1'b0,x168})+$signed({1'b0,x353})+$signed({1'b0,x297})+$signed(-{1'b0,x224})+$signed(-{1'b0,x104})+$signed(-{2'b0,x105}<<<3'd1)+$signed(sharing70)+$signed(sharing71)-$signed(11'd16);
assign y107=temp_y[107][11] ==1'b1 ? 5'd0 :  
        temp_y[107][9] ==1'b1 ? 5'd31 : 
        temp_y[107][3]==1'b1 ? temp_y[107][8:4]+1'b1 : temp_y[107][8:4];
assign temp_y[108] = 
$signed({3'b0,x168}<<<3'd2)+$signed(-{2'b0,x40}<<<3'd1)+$signed({1'b0,x352})+$signed(-{1'b0,x232})+$signed(-{2'b0,x160}<<<3'd1)+$signed(-{2'b0,x233}<<<3'd1)+$signed(-{2'b0,x97}<<<3'd1)+$signed(-{2'b0,x353}<<<3'd1)+$signed(sharing70)+$signed(-sharing71)-$signed(11'd24);
assign y108=temp_y[108][11] ==1'b1 ? 5'd0 :  
        temp_y[108][9] ==1'b1 ? 5'd31 : 
        temp_y[108][3]==1'b1 ? temp_y[108][8:4]+1'b1 : temp_y[108][8:4];
assign temp_y[109] = 
$signed({2'b0,x296}<<<3'd1)+$signed({1'b0,x232})+$signed(-{1'b0,x32})+$signed({3'b0,x297}<<<3'd2)+$signed(-{1'b0,x352})+$signed(-{1'b0,x225})+$signed(-{1'b0,x361})+$signed(-{1'b0,x33})+$signed(-{1'b0,x104})+$signed(-{1'b0,x224})+$signed(-sharing4)-$signed(11'd32);
assign y109=temp_y[109][11] ==1'b1 ? 5'd0 :  
        temp_y[109][9] ==1'b1 ? 5'd31 : 
        temp_y[109][3]==1'b1 ? temp_y[109][8:4]+1'b1 : temp_y[109][8:4];
assign temp_y[110] = 
$signed(-{1'b0,x96})+$signed({3'b0,x353}<<<3'd2)+$signed(-{2'b0,x297}<<<3'd1)+$signed(-{1'b0,x33})+$signed(-{2'b0,x289}<<<3'd1)+$signed({3'b0,x361}<<<3'd2)+$signed(-{1'b0,x41})+$signed(sharing58)-$signed(11'd0);
assign y110=temp_y[110][11] ==1'b1 ? 5'd0 :  
        temp_y[110][9] ==1'b1 ? 5'd31 : 
        temp_y[110][3]==1'b1 ? temp_y[110][8:4]+1'b1 : temp_y[110][8:4];
assign temp_y[111] = 
$signed(-{2'b0,x288}<<<3'd1)+$signed({1'b0,x224})+$signed(-{1'b0,x160})+$signed({3'b0,x105}<<<3'd2)+$signed({2'b0,x353}<<<3'd1)+$signed({1'b0,x289})+$signed(-{3'b0,x361}<<<3'd2)+$signed(-{1'b0,x225})+$signed(-{1'b0,x360})+$signed(-sharing83)-$signed(11'd0);
assign y111=temp_y[111][11] ==1'b1 ? 5'd0 :  
        temp_y[111][9] ==1'b1 ? 5'd31 : 
        temp_y[111][3]==1'b1 ? temp_y[111][8:4]+1'b1 : temp_y[111][8:4];
assign temp_y[112] = 
$signed(-{3'b0,x40}<<<3'd2)+$signed(-{2'b0,x224}<<<3'd1)+$signed(-{1'b0,x296})+$signed({1'b0,x360})+$signed(-{1'b0,x168})+$signed({2'b0,x225}<<<3'd1)+$signed(-{2'b0,x41}<<<3'd1)+$signed(-{2'b0,x169}<<<3'd1)+$signed(-{2'b0,x32}<<<3'd1)+$signed({1'b0,x96})+$signed(sharing15)+$signed(11'd40);
assign y112=temp_y[112][11] ==1'b1 ? 5'd0 :  
        temp_y[112][9] ==1'b1 ? 5'd31 : 
        temp_y[112][3]==1'b1 ? temp_y[112][8:4]+1'b1 : temp_y[112][8:4];
assign temp_y[113] = 
$signed(-{2'b0,x40}<<<3'd1)+$signed({1'b0,x224})+$signed({4'b0,x41}<<<3'd3)+$signed(-{2'b0,x32}<<<3'd1)+$signed(-{2'b0,x233}<<<3'd1)+$signed(-{1'b0,x225})+$signed(-{1'b0,x361})+$signed({1'b0,x96})+$signed(-sharing15)-$signed(11'd8);
assign y113=temp_y[113][11] ==1'b1 ? 5'd0 :  
        temp_y[113][9] ==1'b1 ? 5'd31 : 
        temp_y[113][3]==1'b1 ? temp_y[113][8:4]+1'b1 : temp_y[113][8:4];
assign temp_y[114] = 
$signed({3'b0,x352}<<<3'd2)+$signed(-{2'b0,x32}<<<3'd1)+$signed(-{1'b0,x168})+$signed({3'b0,x360}<<<3'd2)+$signed(-{1'b0,x40})+$signed({2'b0,x161}<<<3'd1)+$signed({2'b0,x41}<<<3'd1)+$signed({1'b0,x169})+$signed(-{2'b0,x232}<<<3'd1)+$signed(-{2'b0,x297}<<<3'd1)+$signed(-{1'b0,x97})+$signed(-{1'b0,x105})+$signed(-{1'b0,x289})+$signed(-{1'b0,x224})+$signed(-{1'b0,x296})+$signed(-{1'b0,x104})+$signed(sharing4)-$signed(11'd16);
assign y114=temp_y[114][11] ==1'b1 ? 5'd0 :  
        temp_y[114][9] ==1'b1 ? 5'd31 : 
        temp_y[114][3]==1'b1 ? temp_y[114][8:4]+1'b1 : temp_y[114][8:4];
assign temp_y[115] = 
$signed(-{4'b0,x296}<<<3'd3)+$signed(-{3'b0,x224}<<<3'd2)+$signed(-{3'b0,x288}<<<3'd2)+$signed(-{1'b0,x232})+$signed(-{4'b0,x289}<<<3'd3)+$signed(-{4'b0,x233}<<<3'd3)+$signed(-{1'b0,x360})+$signed({1'b0,x41})+$signed(-{1'b0,x105})+$signed(-{1'b0,x351})+$signed(-{1'b0,x225})+$signed(-{1'b0,x359})+$signed(sharing83)+$signed(11'd24);
assign y115=temp_y[115][11] ==1'b1 ? 5'd0 :  
        temp_y[115][9] ==1'b1 ? 5'd31 : 
        temp_y[115][3]==1'b1 ? temp_y[115][8:4]+1'b1 : temp_y[115][8:4];
assign temp_y[116] = 
$signed({3'b0,x232}<<<3'd2)+$signed(-{2'b0,x296}<<<3'd1)+$signed({2'b0,x160}<<<3'd1)+$signed({1'b0,x360})+$signed({2'b0,x352}<<<3'd1)+$signed(-{1'b0,x40})+$signed(-{1'b0,x353})+$signed(-{3'b0,x161}<<<3'd2)+$signed(-{2'b0,x97}<<<3'd1)+$signed(-{3'b0,x169}<<<3'd2)+$signed(-{1'b0,x289})+$signed({1'b0,x41})+$signed({1'b0,x96})+$signed(sharing58)+$signed(11'd16);
assign y116=temp_y[116][11] ==1'b1 ? 5'd0 :  
        temp_y[116][9] ==1'b1 ? 5'd31 : 
        temp_y[116][3]==1'b1 ? temp_y[116][8:4]+1'b1 : temp_y[116][8:4];
assign temp_y[117] = 
$signed(-{3'b0,x362}<<<3'd2)+$signed({2'b0,x298}<<<3'd1)+$signed(-{1'b0,x106})+$signed(-{2'b0,x354}<<<3'd1)+$signed({1'b0,x170})+$signed({2'b0,x291}<<<3'd1)+$signed({1'b0,x299})+$signed(-{1'b0,x107})+$signed(-{1'b0,x163})+$signed(-{3'b0,x363}<<<3'd2)+$signed(sharing43)+$signed(11'd32);
assign y117=temp_y[117][11] ==1'b1 ? 5'd0 :  
        temp_y[117][9] ==1'b1 ? 5'd31 : 
        temp_y[117][3]==1'b1 ? temp_y[117][8:4]+1'b1 : temp_y[117][8:4];
assign temp_y[118] = 
$signed({2'b0,x106}<<<3'd1)+$signed({2'b0,x362}<<<3'd1)+$signed({2'b0,x234}<<<3'd1)+$signed({1'b0,x98})+$signed({1'b0,x34})+$signed(-{1'b0,x35})+$signed(-{1'b0,x298})+$signed(-{2'b0,x235}<<<3'd1)+$signed(-{1'b0,x291})+$signed(-{1'b0,x170})+$signed({3'b0,x363}<<<3'd2)+$signed(sharing43)-$signed(11'd0);
assign y118=temp_y[118][11] ==1'b1 ? 5'd0 :  
        temp_y[118][9] ==1'b1 ? 5'd31 : 
        temp_y[118][3]==1'b1 ? temp_y[118][8:4]+1'b1 : temp_y[118][8:4];
assign temp_y[119] = 
$signed(-{3'b0,x290}<<<3'd2)+$signed(-{2'b0,x106}<<<3'd1)+$signed({2'b0,x234}<<<3'd1)+$signed({1'b0,x162})+$signed({1'b0,x226})+$signed(-{2'b0,x98}<<<3'd1)+$signed(-{4'b0,x291}<<<3'd3)+$signed(-{3'b0,x298}<<<3'd2)+$signed(-{3'b0,x299}<<<3'd2)+$signed(-{1'b0,x235})+$signed(-{1'b0,x171})+$signed(-{3'b0,x362}<<<3'd2)+$signed(-{2'b0,x354}<<<3'd1)+$signed(11'd40);
assign y119=temp_y[119][11] ==1'b1 ? 5'd0 :  
        temp_y[119][9] ==1'b1 ? 5'd31 : 
        temp_y[119][3]==1'b1 ? temp_y[119][8:4]+1'b1 : temp_y[119][8:4];
assign temp_y[120] = 
$signed({2'b0,x354}<<<3'd1)+$signed(-{1'b0,x98})+$signed({1'b0,x42})+$signed({1'b0,x290})+$signed({1'b0,x170})+$signed({1'b0,x355})+$signed({1'b0,x299})+$signed(-{1'b0,x226})+$signed(-{1'b0,x106})+$signed(-{2'b0,x107}<<<3'd1)+$signed(sharing87)+$signed(sharing88)-$signed(11'd16);
assign y120=temp_y[120][11] ==1'b1 ? 5'd0 :  
        temp_y[120][9] ==1'b1 ? 5'd31 : 
        temp_y[120][3]==1'b1 ? temp_y[120][8:4]+1'b1 : temp_y[120][8:4];
assign temp_y[121] = 
$signed({3'b0,x170}<<<3'd2)+$signed(-{2'b0,x42}<<<3'd1)+$signed({1'b0,x354})+$signed(-{1'b0,x234})+$signed(-{2'b0,x162}<<<3'd1)+$signed(-{2'b0,x235}<<<3'd1)+$signed(-{2'b0,x99}<<<3'd1)+$signed(-{2'b0,x355}<<<3'd1)+$signed(sharing87)+$signed(-sharing88)-$signed(11'd24);
assign y121=temp_y[121][11] ==1'b1 ? 5'd0 :  
        temp_y[121][9] ==1'b1 ? 5'd31 : 
        temp_y[121][3]==1'b1 ? temp_y[121][8:4]+1'b1 : temp_y[121][8:4];
assign temp_y[122] = 
$signed({2'b0,x298}<<<3'd1)+$signed(-{1'b0,x34})+$signed({1'b0,x234})+$signed(-{1'b0,x354})+$signed({3'b0,x299}<<<3'd2)+$signed(-{1'b0,x227})+$signed(-{1'b0,x363})+$signed(-{1'b0,x35})+$signed(-{1'b0,x106})+$signed(-{1'b0,x226})+$signed(sharing28)-$signed(11'd32);
assign y122=temp_y[122][11] ==1'b1 ? 5'd0 :  
        temp_y[122][9] ==1'b1 ? 5'd31 : 
        temp_y[122][3]==1'b1 ? temp_y[122][8:4]+1'b1 : temp_y[122][8:4];
assign temp_y[123] = 
$signed(-{1'b0,x98})+$signed({3'b0,x363}<<<3'd2)+$signed(-{2'b0,x291}<<<3'd1)+$signed({3'b0,x355}<<<3'd2)+$signed(-{2'b0,x299}<<<3'd1)+$signed(-{1'b0,x35})+$signed(-{1'b0,x43})+$signed(sharing53)-$signed(11'd0);
assign y123=temp_y[123][11] ==1'b1 ? 5'd0 :  
        temp_y[123][9] ==1'b1 ? 5'd31 : 
        temp_y[123][3]==1'b1 ? temp_y[123][8:4]+1'b1 : temp_y[123][8:4];
assign temp_y[124] = 
$signed(-{2'b0,x290}<<<3'd1)+$signed({1'b0,x226})+$signed(-{1'b0,x162})+$signed(-{3'b0,x363}<<<3'd2)+$signed({3'b0,x107}<<<3'd2)+$signed({2'b0,x355}<<<3'd1)+$signed({1'b0,x291})+$signed(-{1'b0,x227})+$signed(-{1'b0,x362})+$signed(-sharing111)-$signed(11'd0);
assign y124=temp_y[124][11] ==1'b1 ? 5'd0 :  
        temp_y[124][9] ==1'b1 ? 5'd31 : 
        temp_y[124][3]==1'b1 ? temp_y[124][8:4]+1'b1 : temp_y[124][8:4];
assign temp_y[125] = 
$signed(-{3'b0,x42}<<<3'd2)+$signed(-{2'b0,x226}<<<3'd1)+$signed(-{1'b0,x298})+$signed({1'b0,x362})+$signed(-{1'b0,x170})+$signed({2'b0,x227}<<<3'd1)+$signed(-{2'b0,x43}<<<3'd1)+$signed(-{2'b0,x171}<<<3'd1)+$signed(-{2'b0,x34}<<<3'd1)+$signed({1'b0,x98})+$signed(sharing29)+$signed(11'd40);
assign y125=temp_y[125][11] ==1'b1 ? 5'd0 :  
        temp_y[125][9] ==1'b1 ? 5'd31 : 
        temp_y[125][3]==1'b1 ? temp_y[125][8:4]+1'b1 : temp_y[125][8:4];
assign temp_y[126] = 
$signed(-{2'b0,x42}<<<3'd1)+$signed({1'b0,x226})+$signed({4'b0,x43}<<<3'd3)+$signed(-{2'b0,x34}<<<3'd1)+$signed(-{2'b0,x235}<<<3'd1)+$signed(-{1'b0,x227})+$signed(-{1'b0,x363})+$signed({1'b0,x98})+$signed(-sharing29)-$signed(11'd8);
assign y126=temp_y[126][11] ==1'b1 ? 5'd0 :  
        temp_y[126][9] ==1'b1 ? 5'd31 : 
        temp_y[126][3]==1'b1 ? temp_y[126][8:4]+1'b1 : temp_y[126][8:4];
assign temp_y[127] = 
$signed(-{1'b0,x106})+$signed({3'b0,x354}<<<3'd2)+$signed(-{2'b0,x34}<<<3'd1)+$signed(-{1'b0,x170})+$signed({3'b0,x362}<<<3'd2)+$signed(-{1'b0,x42})+$signed({2'b0,x163}<<<3'd1)+$signed({2'b0,x43}<<<3'd1)+$signed({1'b0,x171})+$signed(-{2'b0,x234}<<<3'd1)+$signed(-{2'b0,x299}<<<3'd1)+$signed(-{1'b0,x99})+$signed(-{1'b0,x107})+$signed(-{1'b0,x291})+$signed(-{1'b0,x226})+$signed(-{1'b0,x298})+$signed(-sharing28)-$signed(11'd16);
assign y127=temp_y[127][11] ==1'b1 ? 5'd0 :  
        temp_y[127][9] ==1'b1 ? 5'd31 : 
        temp_y[127][3]==1'b1 ? temp_y[127][8:4]+1'b1 : temp_y[127][8:4];
assign temp_y[128] = 
$signed(-{1'b0,x353})+$signed(-{4'b0,x298}<<<3'd3)+$signed(-{3'b0,x226}<<<3'd2)+$signed(-{3'b0,x290}<<<3'd2)+$signed(-{1'b0,x361})+$signed(-{4'b0,x291}<<<3'd3)+$signed(-{1'b0,x234})+$signed(-{4'b0,x235}<<<3'd3)+$signed({1'b0,x43})+$signed(-{1'b0,x107})+$signed(-{1'b0,x227})+$signed(-{1'b0,x362})+$signed(sharing111)+$signed(11'd24);
assign y128=temp_y[128][11] ==1'b1 ? 5'd0 :  
        temp_y[128][9] ==1'b1 ? 5'd31 : 
        temp_y[128][3]==1'b1 ? temp_y[128][8:4]+1'b1 : temp_y[128][8:4];
assign temp_y[129] = 
$signed({1'b0,x98})+$signed({3'b0,x234}<<<3'd2)+$signed({2'b0,x162}<<<3'd1)+$signed({1'b0,x362})+$signed({2'b0,x354}<<<3'd1)+$signed(-{3'b0,x171}<<<3'd2)+$signed(-{2'b0,x298}<<<3'd1)+$signed(-{1'b0,x355})+$signed(-{1'b0,x42})+$signed(-{3'b0,x163}<<<3'd2)+$signed(-{2'b0,x99}<<<3'd1)+$signed(-{1'b0,x291})+$signed({1'b0,x43})+$signed(sharing53)+$signed(11'd16);
assign y129=temp_y[129][11] ==1'b1 ? 5'd0 :  
        temp_y[129][9] ==1'b1 ? 5'd31 : 
        temp_y[129][3]==1'b1 ? temp_y[129][8:4]+1'b1 : temp_y[129][8:4];
assign temp_y[130] = 
$signed(-{1'b0,x109})+$signed(-{3'b0,x364}<<<3'd2)+$signed({2'b0,x300}<<<3'd1)+$signed(-{2'b0,x356}<<<3'd1)+$signed(-{1'b0,x108})+$signed({1'b0,x172})+$signed({2'b0,x293}<<<3'd1)+$signed(-{1'b0,x165})+$signed(-{3'b0,x365}<<<3'd2)+$signed({1'b0,x301})+$signed(sharing47)+$signed(11'd32);
assign y130=temp_y[130][11] ==1'b1 ? 5'd0 :  
        temp_y[130][9] ==1'b1 ? 5'd31 : 
        temp_y[130][3]==1'b1 ? temp_y[130][8:4]+1'b1 : temp_y[130][8:4];
assign temp_y[131] = 
$signed({2'b0,x236}<<<3'd1)+$signed({2'b0,x108}<<<3'd1)+$signed({2'b0,x364}<<<3'd1)+$signed({1'b0,x36})+$signed({1'b0,x100})+$signed(-{1'b0,x37})+$signed(-{1'b0,x300})+$signed(-{2'b0,x237}<<<3'd1)+$signed(-{1'b0,x293})+$signed(-{1'b0,x172})+$signed({3'b0,x365}<<<3'd2)+$signed(sharing47)-$signed(11'd0);
assign y131=temp_y[131][11] ==1'b1 ? 5'd0 :  
        temp_y[131][9] ==1'b1 ? 5'd31 : 
        temp_y[131][3]==1'b1 ? temp_y[131][8:4]+1'b1 : temp_y[131][8:4];
assign temp_y[132] = 
$signed(-{1'b0,x173})+$signed(-{3'b0,x364}<<<3'd2)+$signed({2'b0,x236}<<<3'd1)+$signed(-{2'b0,x356}<<<3'd1)+$signed({1'b0,x164})+$signed(-{3'b0,x292}<<<3'd2)+$signed({1'b0,x228})+$signed(-{2'b0,x108}<<<3'd1)+$signed(-{2'b0,x100}<<<3'd1)+$signed(-{4'b0,x293}<<<3'd3)+$signed(-{3'b0,x300}<<<3'd2)+$signed(-{3'b0,x301}<<<3'd2)+$signed(-{1'b0,x237})+$signed(11'd40);
assign y132=temp_y[132][11] ==1'b1 ? 5'd0 :  
        temp_y[132][9] ==1'b1 ? 5'd31 : 
        temp_y[132][3]==1'b1 ? temp_y[132][8:4]+1'b1 : temp_y[132][8:4];
assign temp_y[133] = 
$signed({2'b0,x356}<<<3'd1)+$signed(-{1'b0,x100})+$signed({1'b0,x44})+$signed({1'b0,x292})+$signed({1'b0,x172})+$signed({1'b0,x357})+$signed(-{1'b0,x228})+$signed({1'b0,x301})+$signed(-{1'b0,x108})+$signed(-{2'b0,x109}<<<3'd1)+$signed(sharing65)+$signed(sharing66)-$signed(11'd16);
assign y133=temp_y[133][11] ==1'b1 ? 5'd0 :  
        temp_y[133][9] ==1'b1 ? 5'd31 : 
        temp_y[133][3]==1'b1 ? temp_y[133][8:4]+1'b1 : temp_y[133][8:4];
assign temp_y[134] = 
$signed({3'b0,x172}<<<3'd2)+$signed(-{2'b0,x44}<<<3'd1)+$signed({1'b0,x356})+$signed(-{1'b0,x236})+$signed(-{2'b0,x164}<<<3'd1)+$signed(-{2'b0,x237}<<<3'd1)+$signed(-{2'b0,x101}<<<3'd1)+$signed(-{2'b0,x357}<<<3'd1)+$signed(sharing65)+$signed(-sharing66)-$signed(11'd24);
assign y134=temp_y[134][11] ==1'b1 ? 5'd0 :  
        temp_y[134][9] ==1'b1 ? 5'd31 : 
        temp_y[134][3]==1'b1 ? temp_y[134][8:4]+1'b1 : temp_y[134][8:4];
assign temp_y[135] = 
$signed(-{1'b0,x365})+$signed({2'b0,x300}<<<3'd1)+$signed({1'b0,x236})+$signed(-{1'b0,x36})+$signed({3'b0,x301}<<<3'd2)+$signed(-{1'b0,x356})+$signed(-{1'b0,x229})+$signed(-{1'b0,x37})+$signed(-{1'b0,x108})+$signed(-{1'b0,x228})+$signed(-sharing32)-$signed(11'd32);
assign y135=temp_y[135][11] ==1'b1 ? 5'd0 :  
        temp_y[135][9] ==1'b1 ? 5'd31 : 
        temp_y[135][3]==1'b1 ? temp_y[135][8:4]+1'b1 : temp_y[135][8:4];
assign temp_y[136] = 
$signed(-{1'b0,x100})+$signed({3'b0,x357}<<<3'd2)+$signed(-{2'b0,x301}<<<3'd1)+$signed(-{1'b0,x37})+$signed(-{2'b0,x293}<<<3'd1)+$signed({3'b0,x365}<<<3'd2)+$signed(-{1'b0,x45})+$signed(sharing50)-$signed(11'd0);
assign y136=temp_y[136][11] ==1'b1 ? 5'd0 :  
        temp_y[136][9] ==1'b1 ? 5'd31 : 
        temp_y[136][3]==1'b1 ? temp_y[136][8:4]+1'b1 : temp_y[136][8:4];
assign temp_y[137] = 
$signed(-{1'b0,x229})+$signed(-{2'b0,x292}<<<3'd1)+$signed({1'b0,x228})+$signed(-{1'b0,x164})+$signed({3'b0,x109}<<<3'd2)+$signed({2'b0,x357}<<<3'd1)+$signed({1'b0,x293})+$signed(-{3'b0,x365}<<<3'd2)+$signed(-{1'b0,x364})+$signed(sharing104)-$signed(11'd0);
assign y137=temp_y[137][11] ==1'b1 ? 5'd0 :  
        temp_y[137][9] ==1'b1 ? 5'd31 : 
        temp_y[137][3]==1'b1 ? temp_y[137][8:4]+1'b1 : temp_y[137][8:4];
assign temp_y[138] = 
$signed(-{3'b0,x44}<<<3'd2)+$signed(-{2'b0,x228}<<<3'd1)+$signed(-{1'b0,x300})+$signed({1'b0,x364})+$signed(-{1'b0,x172})+$signed({2'b0,x229}<<<3'd1)+$signed(-{2'b0,x45}<<<3'd1)+$signed(-{2'b0,x173}<<<3'd1)+$signed(-{2'b0,x36}<<<3'd1)+$signed({1'b0,x100})+$signed(sharing13)+$signed(11'd40);
assign y138=temp_y[138][11] ==1'b1 ? 5'd0 :  
        temp_y[138][9] ==1'b1 ? 5'd31 : 
        temp_y[138][3]==1'b1 ? temp_y[138][8:4]+1'b1 : temp_y[138][8:4];
assign temp_y[139] = 
$signed(-{1'b0,x229})+$signed(-{2'b0,x44}<<<3'd1)+$signed({1'b0,x228})+$signed({4'b0,x45}<<<3'd3)+$signed(-{2'b0,x36}<<<3'd1)+$signed(-{2'b0,x237}<<<3'd1)+$signed(-{1'b0,x365})+$signed({1'b0,x100})+$signed(-sharing13)-$signed(11'd8);
assign y139=temp_y[139][11] ==1'b1 ? 5'd0 :  
        temp_y[139][9] ==1'b1 ? 5'd31 : 
        temp_y[139][3]==1'b1 ? temp_y[139][8:4]+1'b1 : temp_y[139][8:4];
assign temp_y[140] = 
$signed(-{1'b0,x101})+$signed(-{1'b0,x109})+$signed({1'b0,x173})+$signed(-{1'b0,x228})+$signed({3'b0,x356}<<<3'd2)+$signed({3'b0,x364}<<<3'd2)+$signed(-{2'b0,x36}<<<3'd1)+$signed(-{1'b0,x44})+$signed(-{1'b0,x172})+$signed({2'b0,x165}<<<3'd1)+$signed(-{1'b0,x293})+$signed({2'b0,x45}<<<3'd1)+$signed(-{2'b0,x236}<<<3'd1)+$signed(-{1'b0,x300})+$signed(-{2'b0,x301}<<<3'd1)+$signed(-{1'b0,x108})+$signed(sharing32)-$signed(11'd16);
assign y140=temp_y[140][11] ==1'b1 ? 5'd0 :  
        temp_y[140][9] ==1'b1 ? 5'd31 : 
        temp_y[140][3]==1'b1 ? temp_y[140][8:4]+1'b1 : temp_y[140][8:4];
assign temp_y[141] = 
$signed(-{1'b0,x355})+$signed(-{1'b0,x363})+$signed(-{3'b0,x228}<<<3'd2)+$signed(-{3'b0,x292}<<<3'd2)+$signed(-{4'b0,x300}<<<3'd3)+$signed(-{4'b0,x293}<<<3'd3)+$signed(-{1'b0,x236})+$signed(-{4'b0,x237}<<<3'd3)+$signed(-{1'b0,x109})+$signed(-{1'b0,x229})+$signed({1'b0,x45})+$signed(-{1'b0,x364})+$signed(-sharing104)+$signed(11'd24);
assign y141=temp_y[141][11] ==1'b1 ? 5'd0 :  
        temp_y[141][9] ==1'b1 ? 5'd31 : 
        temp_y[141][3]==1'b1 ? temp_y[141][8:4]+1'b1 : temp_y[141][8:4];
assign temp_y[142] = 
$signed(-{1'b0,x293})+$signed({3'b0,x236}<<<3'd2)+$signed({2'b0,x164}<<<3'd1)+$signed({1'b0,x364})+$signed({2'b0,x356}<<<3'd1)+$signed(-{2'b0,x300}<<<3'd1)+$signed(-{1'b0,x44})+$signed(-{1'b0,x357})+$signed(-{3'b0,x165}<<<3'd2)+$signed(-{2'b0,x101}<<<3'd1)+$signed(-{3'b0,x173}<<<3'd2)+$signed({1'b0,x100})+$signed({1'b0,x45})+$signed(sharing50)+$signed(11'd16);
assign y142=temp_y[142][11] ==1'b1 ? 5'd0 :  
        temp_y[142][9] ==1'b1 ? 5'd31 : 
        temp_y[142][3]==1'b1 ? temp_y[142][8:4]+1'b1 : temp_y[142][8:4];
assign temp_y[143] = 
$signed({1'b0,x303})+$signed({2'b0,x302}<<<3'd1)+$signed(-{1'b0,x111})+$signed(-{3'b0,x367}<<<3'd2)+$signed(-{3'b0,x366}<<<3'd2)+$signed(-{2'b0,x358}<<<3'd1)+$signed(-{1'b0,x110})+$signed({1'b0,x174})+$signed({2'b0,x295}<<<3'd1)+$signed(-{1'b0,x167})+$signed(sharing33)+$signed(11'd32);
assign y143=temp_y[143][11] ==1'b1 ? 5'd0 :  
        temp_y[143][9] ==1'b1 ? 5'd31 : 
        temp_y[143][3]==1'b1 ? temp_y[143][8:4]+1'b1 : temp_y[143][8:4];
assign temp_y[144] = 
$signed({2'b0,x238}<<<3'd1)+$signed(-{1'b0,x295})+$signed(-{1'b0,x302})+$signed({2'b0,x366}<<<3'd1)+$signed({3'b0,x367}<<<3'd2)+$signed({1'b0,x102})+$signed({2'b0,x110}<<<3'd1)+$signed({1'b0,x38})+$signed(-{1'b0,x174})+$signed(-{2'b0,x239}<<<3'd1)+$signed(-{1'b0,x39})+$signed(sharing33)-$signed(11'd0);
assign y144=temp_y[144][11] ==1'b1 ? 5'd0 :  
        temp_y[144][9] ==1'b1 ? 5'd31 : 
        temp_y[144][3]==1'b1 ? temp_y[144][8:4]+1'b1 : temp_y[144][8:4];
assign temp_y[145] = 
$signed({2'b0,x238}<<<3'd1)+$signed(-{3'b0,x302}<<<3'd2)+$signed(-{3'b0,x366}<<<3'd2)+$signed(-{2'b0,x358}<<<3'd1)+$signed(-{2'b0,x110}<<<3'd1)+$signed(-{4'b0,x295}<<<3'd3)+$signed(-{1'b0,x175})+$signed(-{3'b0,x294}<<<3'd2)+$signed(-{2'b0,x102}<<<3'd1)+$signed({1'b0,x230})+$signed({1'b0,x166})+$signed(-{3'b0,x303}<<<3'd2)+$signed(-{1'b0,x239})+$signed(11'd40);
assign y145=temp_y[145][11] ==1'b1 ? 5'd0 :  
        temp_y[145][9] ==1'b1 ? 5'd31 : 
        temp_y[145][3]==1'b1 ? temp_y[145][8:4]+1'b1 : temp_y[145][8:4];
assign temp_y[146] = 
$signed(-{1'b0,x230})+$signed({1'b0,x359})+$signed({1'b0,x294})+$signed({1'b0,x46})+$signed(-{1'b0,x102})+$signed({2'b0,x358}<<<3'd1)+$signed(-{1'b0,x110})+$signed({1'b0,x174})+$signed(-{2'b0,x111}<<<3'd1)+$signed({1'b0,x303})+$signed(sharing84)+$signed(sharing85)-$signed(11'd16);
assign y146=temp_y[146][11] ==1'b1 ? 5'd0 :  
        temp_y[146][9] ==1'b1 ? 5'd31 : 
        temp_y[146][3]==1'b1 ? temp_y[146][8:4]+1'b1 : temp_y[146][8:4];
assign temp_y[147] = 
$signed(-{2'b0,x103}<<<3'd1)+$signed(-{2'b0,x359}<<<3'd1)+$signed({1'b0,x358})+$signed(-{2'b0,x166}<<<3'd1)+$signed({3'b0,x174}<<<3'd2)+$signed(-{2'b0,x46}<<<3'd1)+$signed(-{1'b0,x238})+$signed(-{2'b0,x239}<<<3'd1)+$signed(sharing84)+$signed(-sharing85)-$signed(11'd24);
assign y147=temp_y[147][11] ==1'b1 ? 5'd0 :  
        temp_y[147][9] ==1'b1 ? 5'd31 : 
        temp_y[147][3]==1'b1 ? temp_y[147][8:4]+1'b1 : temp_y[147][8:4];
assign temp_y[148] = 
$signed(-{1'b0,x39})+$signed(-{1'b0,x230})+$signed({1'b0,x238})+$signed(-{1'b0,x367})+$signed(-{1'b0,x358})+$signed(-{1'b0,x110})+$signed({2'b0,x302}<<<3'd1)+$signed(-{1'b0,x38})+$signed({3'b0,x303}<<<3'd2)+$signed(-{1'b0,x231})+$signed(-sharing9)-$signed(11'd32);
assign y148=temp_y[148][11] ==1'b1 ? 5'd0 :  
        temp_y[148][9] ==1'b1 ? 5'd31 : 
        temp_y[148][3]==1'b1 ? temp_y[148][8:4]+1'b1 : temp_y[148][8:4];
assign temp_y[149] = 
$signed(-{1'b0,x47})+$signed({3'b0,x359}<<<3'd2)+$signed(-{1'b0,x102})+$signed(-{2'b0,x303}<<<3'd1)+$signed({3'b0,x367}<<<3'd2)+$signed(-{2'b0,x295}<<<3'd1)+$signed(-{1'b0,x39})+$signed(sharing51)-$signed(11'd0);
assign y149=temp_y[149][11] ==1'b1 ? 5'd0 :  
        temp_y[149][9] ==1'b1 ? 5'd31 : 
        temp_y[149][3]==1'b1 ? temp_y[149][8:4]+1'b1 : temp_y[149][8:4];
assign temp_y[150] = 
$signed({1'b0,x295})+$signed(-{1'b0,x366})+$signed(-{1'b0,x231})+$signed(-{2'b0,x294}<<<3'd1)+$signed({1'b0,x230})+$signed(-{1'b0,x166})+$signed(-{3'b0,x367}<<<3'd2)+$signed({2'b0,x359}<<<3'd1)+$signed({3'b0,x111}<<<3'd2)+$signed(-sharing108)-$signed(11'd0);
assign y150=temp_y[150][11] ==1'b1 ? 5'd0 :  
        temp_y[150][9] ==1'b1 ? 5'd31 : 
        temp_y[150][3]==1'b1 ? temp_y[150][8:4]+1'b1 : temp_y[150][8:4];
assign temp_y[151] = 
$signed(-{2'b0,x38}<<<3'd1)+$signed({2'b0,x231}<<<3'd1)+$signed({1'b0,x102})+$signed({1'b0,x366})+$signed(-{3'b0,x46}<<<3'd2)+$signed(-{2'b0,x230}<<<3'd1)+$signed(-{1'b0,x302})+$signed(-{2'b0,x47}<<<3'd1)+$signed(-{1'b0,x174})+$signed(-{2'b0,x175}<<<3'd1)+$signed(-sharing18)+$signed(11'd40);
assign y151=temp_y[151][11] ==1'b1 ? 5'd0 :  
        temp_y[151][9] ==1'b1 ? 5'd31 : 
        temp_y[151][3]==1'b1 ? temp_y[151][8:4]+1'b1 : temp_y[151][8:4];
assign temp_y[152] = 
$signed(-{2'b0,x38}<<<3'd1)+$signed(-{1'b0,x367})+$signed({1'b0,x102})+$signed(-{2'b0,x46}<<<3'd1)+$signed({1'b0,x230})+$signed({4'b0,x47}<<<3'd3)+$signed(-{2'b0,x239}<<<3'd1)+$signed(-{1'b0,x231})+$signed(sharing18)-$signed(11'd8);
assign y152=temp_y[152][11] ==1'b1 ? 5'd0 :  
        temp_y[152][9] ==1'b1 ? 5'd31 : 
        temp_y[152][3]==1'b1 ? temp_y[152][8:4]+1'b1 : temp_y[152][8:4];
assign temp_y[153] = 
$signed(-{1'b0,x295})+$signed(-{1'b0,x230})+$signed(-{2'b0,x38}<<<3'd1)+$signed(-{1'b0,x111})+$signed({3'b0,x366}<<<3'd2)+$signed({2'b0,x167}<<<3'd1)+$signed(-{1'b0,x46})+$signed({1'b0,x175})+$signed(-{1'b0,x110})+$signed({3'b0,x358}<<<3'd2)+$signed(-{2'b0,x238}<<<3'd1)+$signed(-{1'b0,x302})+$signed({2'b0,x47}<<<3'd1)+$signed(-{1'b0,x174})+$signed(-{2'b0,x303}<<<3'd1)+$signed(-{1'b0,x103})+$signed(sharing9)-$signed(11'd16);
assign y153=temp_y[153][11] ==1'b1 ? 5'd0 :  
        temp_y[153][9] ==1'b1 ? 5'd31 : 
        temp_y[153][3]==1'b1 ? temp_y[153][8:4]+1'b1 : temp_y[153][8:4];
assign temp_y[154] = 
$signed(-{1'b0,x357})+$signed({1'b0,x47})+$signed(-{4'b0,x239}<<<3'd3)+$signed(-{1'b0,x366})+$signed(-{1'b0,x365})+$signed(-{4'b0,x302}<<<3'd3)+$signed(-{3'b0,x294}<<<3'd2)+$signed(-{3'b0,x230}<<<3'd2)+$signed(-{1'b0,x238})+$signed(-{4'b0,x295}<<<3'd3)+$signed(-{1'b0,x231})+$signed(-{1'b0,x111})+$signed(sharing108)+$signed(11'd24);
assign y154=temp_y[154][11] ==1'b1 ? 5'd0 :  
        temp_y[154][9] ==1'b1 ? 5'd31 : 
        temp_y[154][3]==1'b1 ? temp_y[154][8:4]+1'b1 : temp_y[154][8:4];
assign temp_y[155] = 
$signed({1'b0,x47})+$signed(-{3'b0,x175}<<<3'd2)+$signed(-{2'b0,x302}<<<3'd1)+$signed(-{1'b0,x359})+$signed({1'b0,x102})+$signed({1'b0,x366})+$signed({2'b0,x166}<<<3'd1)+$signed({3'b0,x238}<<<3'd2)+$signed({2'b0,x358}<<<3'd1)+$signed(-{1'b0,x46})+$signed(-{3'b0,x167}<<<3'd2)+$signed(-{2'b0,x103}<<<3'd1)+$signed(-{1'b0,x295})+$signed(sharing51)+$signed(11'd16);
assign y155=temp_y[155][11] ==1'b1 ? 5'd0 :  
        temp_y[155][9] ==1'b1 ? 5'd31 : 
        temp_y[155][3]==1'b1 ? temp_y[155][8:4]+1'b1 : temp_y[155][8:4];
assign temp_y[156] = 
$signed(-{3'b0,x376}<<<3'd2)+$signed({2'b0,x312}<<<3'd1)+$signed(-{1'b0,x120})+$signed(-{2'b0,x368}<<<3'd1)+$signed({1'b0,x184})+$signed({2'b0,x305}<<<3'd1)+$signed({1'b0,x313})+$signed(-{1'b0,x177})+$signed(-{1'b0,x121})+$signed(-{3'b0,x377}<<<3'd2)+$signed(sharing42)+$signed(11'd32);
assign y156=temp_y[156][11] ==1'b1 ? 5'd0 :  
        temp_y[156][9] ==1'b1 ? 5'd31 : 
        temp_y[156][3]==1'b1 ? temp_y[156][8:4]+1'b1 : temp_y[156][8:4];
assign temp_y[157] = 
$signed({2'b0,x248}<<<3'd1)+$signed({2'b0,x120}<<<3'd1)+$signed({2'b0,x376}<<<3'd1)+$signed({1'b0,x48})+$signed({1'b0,x112})+$signed(-{1'b0,x305})+$signed(-{1'b0,x312})+$signed(-{2'b0,x249}<<<3'd1)+$signed(-{1'b0,x49})+$signed(-{1'b0,x184})+$signed({3'b0,x377}<<<3'd2)+$signed(sharing42)-$signed(11'd0);
assign y157=temp_y[157][11] ==1'b1 ? 5'd0 :  
        temp_y[157][9] ==1'b1 ? 5'd31 : 
        temp_y[157][3]==1'b1 ? temp_y[157][8:4]+1'b1 : temp_y[157][8:4];
assign temp_y[158] = 
$signed(-{3'b0,x304}<<<3'd2)+$signed({2'b0,x248}<<<3'd1)+$signed({1'b0,x176})+$signed({1'b0,x240})+$signed(-{2'b0,x112}<<<3'd1)+$signed(-{2'b0,x120}<<<3'd1)+$signed(-{4'b0,x305}<<<3'd3)+$signed(-{3'b0,x312}<<<3'd2)+$signed(-{3'b0,x313}<<<3'd2)+$signed(-{1'b0,x249})+$signed(-{1'b0,x185})+$signed(-{3'b0,x376}<<<3'd2)+$signed(-{2'b0,x368}<<<3'd1)+$signed(11'd40);
assign y158=temp_y[158][11] ==1'b1 ? 5'd0 :  
        temp_y[158][9] ==1'b1 ? 5'd31 : 
        temp_y[158][3]==1'b1 ? temp_y[158][8:4]+1'b1 : temp_y[158][8:4];
assign temp_y[159] = 
$signed({2'b0,x368}<<<3'd1)+$signed({1'b0,x304})+$signed({1'b0,x56})+$signed(-{1'b0,x120})+$signed({1'b0,x184})+$signed({1'b0,x369})+$signed({1'b0,x313})+$signed(-{2'b0,x121}<<<3'd1)+$signed(-{1'b0,x112})+$signed(-{1'b0,x240})+$signed(sharing81)+$signed(-sharing82)-$signed(11'd16);
assign y159=temp_y[159][11] ==1'b1 ? 5'd0 :  
        temp_y[159][9] ==1'b1 ? 5'd31 : 
        temp_y[159][3]==1'b1 ? temp_y[159][8:4]+1'b1 : temp_y[159][8:4];
assign temp_y[160] = 
$signed({3'b0,x184}<<<3'd2)+$signed(-{2'b0,x56}<<<3'd1)+$signed(-{2'b0,x176}<<<3'd1)+$signed({1'b0,x368})+$signed(-{1'b0,x248})+$signed(-{2'b0,x249}<<<3'd1)+$signed(-{2'b0,x113}<<<3'd1)+$signed(-{2'b0,x369}<<<3'd1)+$signed(sharing81)+$signed(sharing82)-$signed(11'd24);
assign y160=temp_y[160][11] ==1'b1 ? 5'd0 :  
        temp_y[160][9] ==1'b1 ? 5'd31 : 
        temp_y[160][3]==1'b1 ? temp_y[160][8:4]+1'b1 : temp_y[160][8:4];
assign temp_y[161] = 
$signed({2'b0,x312}<<<3'd1)+$signed(-{1'b0,x368})+$signed({1'b0,x248})+$signed({3'b0,x313}<<<3'd2)+$signed(-{1'b0,x48})+$signed(-{1'b0,x241})+$signed(-{1'b0,x377})+$signed(-{1'b0,x49})+$signed(-{1'b0,x120})+$signed(-{1'b0,x240})+$signed(sharing3)-$signed(11'd32);
assign y161=temp_y[161][11] ==1'b1 ? 5'd0 :  
        temp_y[161][9] ==1'b1 ? 5'd31 : 
        temp_y[161][3]==1'b1 ? temp_y[161][8:4]+1'b1 : temp_y[161][8:4];
assign temp_y[162] = 
$signed(-{1'b0,x112})+$signed({3'b0,x369}<<<3'd2)+$signed(-{2'b0,x313}<<<3'd1)+$signed({3'b0,x377}<<<3'd2)+$signed(-{2'b0,x305}<<<3'd1)+$signed(-{1'b0,x49})+$signed(-{1'b0,x57})+$signed(sharing49)-$signed(11'd0);
assign y162=temp_y[162][11] ==1'b1 ? 5'd0 :  
        temp_y[162][9] ==1'b1 ? 5'd31 : 
        temp_y[162][3]==1'b1 ? temp_y[162][8:4]+1'b1 : temp_y[162][8:4];
assign temp_y[163] = 
$signed(-{2'b0,x304}<<<3'd1)+$signed({1'b0,x240})+$signed(-{1'b0,x176})+$signed({3'b0,x121}<<<3'd2)+$signed({2'b0,x369}<<<3'd1)+$signed({1'b0,x305})+$signed(-{3'b0,x377}<<<3'd2)+$signed(-{1'b0,x241})+$signed(-{1'b0,x376})+$signed(sharing99)-$signed(11'd0);
assign y163=temp_y[163][11] ==1'b1 ? 5'd0 :  
        temp_y[163][9] ==1'b1 ? 5'd31 : 
        temp_y[163][3]==1'b1 ? temp_y[163][8:4]+1'b1 : temp_y[163][8:4];
assign temp_y[164] = 
$signed(-{3'b0,x56}<<<3'd2)+$signed(-{2'b0,x240}<<<3'd1)+$signed({1'b0,x376})+$signed(-{1'b0,x312})+$signed(-{1'b0,x184})+$signed({2'b0,x241}<<<3'd1)+$signed(-{2'b0,x57}<<<3'd1)+$signed(-{2'b0,x185}<<<3'd1)+$signed(-{2'b0,x48}<<<3'd1)+$signed({1'b0,x112})+$signed(sharing1)+$signed(11'd40);
assign y164=temp_y[164][11] ==1'b1 ? 5'd0 :  
        temp_y[164][9] ==1'b1 ? 5'd31 : 
        temp_y[164][3]==1'b1 ? temp_y[164][8:4]+1'b1 : temp_y[164][8:4];
assign temp_y[165] = 
$signed(-{2'b0,x56}<<<3'd1)+$signed({1'b0,x240})+$signed({4'b0,x57}<<<3'd3)+$signed(-{2'b0,x48}<<<3'd1)+$signed(-{2'b0,x249}<<<3'd1)+$signed(-{1'b0,x241})+$signed(-{1'b0,x377})+$signed({1'b0,x112})+$signed(-sharing1)-$signed(11'd8);
assign y165=temp_y[165][11] ==1'b1 ? 5'd0 :  
        temp_y[165][9] ==1'b1 ? 5'd31 : 
        temp_y[165][3]==1'b1 ? temp_y[165][8:4]+1'b1 : temp_y[165][8:4];
assign temp_y[166] = 
$signed({3'b0,x368}<<<3'd2)+$signed(-{2'b0,x48}<<<3'd1)+$signed(-{1'b0,x56})+$signed({3'b0,x376}<<<3'd2)+$signed(-{1'b0,x184})+$signed({2'b0,x177}<<<3'd1)+$signed({1'b0,x185})+$signed({2'b0,x57}<<<3'd1)+$signed(-{2'b0,x248}<<<3'd1)+$signed(-{2'b0,x313}<<<3'd1)+$signed(-{1'b0,x121})+$signed(-{1'b0,x113})+$signed(-{1'b0,x305})+$signed(-{1'b0,x240})+$signed(-{1'b0,x312})+$signed(-{1'b0,x120})+$signed(-sharing3)-$signed(11'd16);
assign y166=temp_y[166][11] ==1'b1 ? 5'd0 :  
        temp_y[166][9] ==1'b1 ? 5'd31 : 
        temp_y[166][3]==1'b1 ? temp_y[166][8:4]+1'b1 : temp_y[166][8:4];
assign temp_y[167] = 
$signed(-{4'b0,x312}<<<3'd3)+$signed(-{3'b0,x240}<<<3'd2)+$signed(-{3'b0,x304}<<<3'd2)+$signed(-{1'b0,x248})+$signed(-{4'b0,x305}<<<3'd3)+$signed(-{4'b0,x249}<<<3'd3)+$signed(-{1'b0,x376})+$signed({1'b0,x57})+$signed(-{1'b0,x121})+$signed(-{1'b0,x367})+$signed(-{1'b0,x241})+$signed(-{1'b0,x375})+$signed(-sharing99)+$signed(11'd24);
assign y167=temp_y[167][11] ==1'b1 ? 5'd0 :  
        temp_y[167][9] ==1'b1 ? 5'd31 : 
        temp_y[167][3]==1'b1 ? temp_y[167][8:4]+1'b1 : temp_y[167][8:4];
assign temp_y[168] = 
$signed({3'b0,x248}<<<3'd2)+$signed({2'b0,x176}<<<3'd1)+$signed({1'b0,x376})+$signed(-{2'b0,x312}<<<3'd1)+$signed({2'b0,x368}<<<3'd1)+$signed(-{1'b0,x56})+$signed(-{1'b0,x369})+$signed(-{3'b0,x185}<<<3'd2)+$signed(-{3'b0,x177}<<<3'd2)+$signed(-{2'b0,x113}<<<3'd1)+$signed(-{1'b0,x305})+$signed({1'b0,x57})+$signed({1'b0,x112})+$signed(sharing49)+$signed(11'd16);
assign y168=temp_y[168][11] ==1'b1 ? 5'd0 :  
        temp_y[168][9] ==1'b1 ? 5'd31 : 
        temp_y[168][3]==1'b1 ? temp_y[168][8:4]+1'b1 : temp_y[168][8:4];
assign temp_y[169] = 
$signed(-{3'b0,x378}<<<3'd2)+$signed({2'b0,x314}<<<3'd1)+$signed(-{1'b0,x122})+$signed(-{2'b0,x370}<<<3'd1)+$signed({1'b0,x186})+$signed({2'b0,x307}<<<3'd1)+$signed({1'b0,x315})+$signed(-{1'b0,x179})+$signed(-{1'b0,x123})+$signed(-{3'b0,x379}<<<3'd2)+$signed(sharing36)+$signed(11'd32);
assign y169=temp_y[169][11] ==1'b1 ? 5'd0 :  
        temp_y[169][9] ==1'b1 ? 5'd31 : 
        temp_y[169][3]==1'b1 ? temp_y[169][8:4]+1'b1 : temp_y[169][8:4];
assign temp_y[170] = 
$signed({2'b0,x250}<<<3'd1)+$signed({2'b0,x122}<<<3'd1)+$signed({1'b0,x114})+$signed({2'b0,x378}<<<3'd1)+$signed({1'b0,x50})+$signed(-{1'b0,x307})+$signed(-{1'b0,x314})+$signed(-{2'b0,x251}<<<3'd1)+$signed(-{1'b0,x51})+$signed(-{1'b0,x186})+$signed({3'b0,x379}<<<3'd2)+$signed(sharing36)-$signed(11'd0);
assign y170=temp_y[170][11] ==1'b1 ? 5'd0 :  
        temp_y[170][9] ==1'b1 ? 5'd31 : 
        temp_y[170][3]==1'b1 ? temp_y[170][8:4]+1'b1 : temp_y[170][8:4];
assign temp_y[171] = 
$signed(-{3'b0,x306}<<<3'd2)+$signed(-{2'b0,x370}<<<3'd1)+$signed({2'b0,x250}<<<3'd1)+$signed({1'b0,x178})+$signed({1'b0,x242})+$signed(-{2'b0,x114}<<<3'd1)+$signed(-{2'b0,x122}<<<3'd1)+$signed(-{4'b0,x307}<<<3'd3)+$signed(-{3'b0,x314}<<<3'd2)+$signed(-{3'b0,x315}<<<3'd2)+$signed(-{1'b0,x251})+$signed(-{1'b0,x187})+$signed(-{3'b0,x378}<<<3'd2)+$signed(11'd40);
assign y171=temp_y[171][11] ==1'b1 ? 5'd0 :  
        temp_y[171][9] ==1'b1 ? 5'd31 : 
        temp_y[171][3]==1'b1 ? temp_y[171][8:4]+1'b1 : temp_y[171][8:4];
assign temp_y[172] = 
$signed({2'b0,x370}<<<3'd1)+$signed({1'b0,x306})+$signed({1'b0,x186})+$signed(-{1'b0,x122})+$signed({1'b0,x58})+$signed({1'b0,x315})+$signed({1'b0,x371})+$signed(-{2'b0,x123}<<<3'd1)+$signed(-{1'b0,x114})+$signed(-{1'b0,x242})+$signed(sharing109)+$signed(sharing110)-$signed(11'd16);
assign y172=temp_y[172][11] ==1'b1 ? 5'd0 :  
        temp_y[172][9] ==1'b1 ? 5'd31 : 
        temp_y[172][3]==1'b1 ? temp_y[172][8:4]+1'b1 : temp_y[172][8:4];
assign temp_y[173] = 
$signed({3'b0,x186}<<<3'd2)+$signed(-{2'b0,x58}<<<3'd1)+$signed(-{2'b0,x178}<<<3'd1)+$signed({1'b0,x370})+$signed(-{1'b0,x250})+$signed(-{2'b0,x251}<<<3'd1)+$signed(-{2'b0,x115}<<<3'd1)+$signed(-{2'b0,x371}<<<3'd1)+$signed(sharing109)+$signed(-sharing110)-$signed(11'd24);
assign y173=temp_y[173][11] ==1'b1 ? 5'd0 :  
        temp_y[173][9] ==1'b1 ? 5'd31 : 
        temp_y[173][3]==1'b1 ? temp_y[173][8:4]+1'b1 : temp_y[173][8:4];
assign temp_y[174] = 
$signed({2'b0,x314}<<<3'd1)+$signed(-{1'b0,x370})+$signed({1'b0,x250})+$signed({3'b0,x315}<<<3'd2)+$signed(-{1'b0,x50})+$signed(-{1'b0,x243})+$signed(-{1'b0,x51})+$signed(-{1'b0,x379})+$signed(-{1'b0,x122})+$signed(-{1'b0,x242})+$signed(-sharing7)-$signed(11'd32);
assign y174=temp_y[174][11] ==1'b1 ? 5'd0 :  
        temp_y[174][9] ==1'b1 ? 5'd31 : 
        temp_y[174][3]==1'b1 ? temp_y[174][8:4]+1'b1 : temp_y[174][8:4];
assign temp_y[175] = 
$signed(-{1'b0,x114})+$signed({3'b0,x379}<<<3'd2)+$signed(-{2'b0,x307}<<<3'd1)+$signed({3'b0,x371}<<<3'd2)+$signed(-{2'b0,x315}<<<3'd1)+$signed(-{1'b0,x51})+$signed(-{1'b0,x59})+$signed(sharing59)-$signed(11'd0);
assign y175=temp_y[175][11] ==1'b1 ? 5'd0 :  
        temp_y[175][9] ==1'b1 ? 5'd31 : 
        temp_y[175][3]==1'b1 ? temp_y[175][8:4]+1'b1 : temp_y[175][8:4];
assign temp_y[176] = 
$signed(-{2'b0,x306}<<<3'd1)+$signed(-{1'b0,x178})+$signed({1'b0,x242})+$signed({3'b0,x123}<<<3'd2)+$signed(-{3'b0,x379}<<<3'd2)+$signed({2'b0,x371}<<<3'd1)+$signed({1'b0,x307})+$signed(-{1'b0,x243})+$signed(-{1'b0,x378})+$signed(sharing80)-$signed(11'd0);
assign y176=temp_y[176][11] ==1'b1 ? 5'd0 :  
        temp_y[176][9] ==1'b1 ? 5'd31 : 
        temp_y[176][3]==1'b1 ? temp_y[176][8:4]+1'b1 : temp_y[176][8:4];
assign temp_y[177] = 
$signed(-{3'b0,x58}<<<3'd2)+$signed(-{2'b0,x242}<<<3'd1)+$signed({1'b0,x378})+$signed(-{1'b0,x314})+$signed(-{1'b0,x186})+$signed({2'b0,x243}<<<3'd1)+$signed(-{2'b0,x59}<<<3'd1)+$signed(-{2'b0,x187}<<<3'd1)+$signed(-{2'b0,x50}<<<3'd1)+$signed({1'b0,x114})+$signed(sharing10)+$signed(11'd40);
assign y177=temp_y[177][11] ==1'b1 ? 5'd0 :  
        temp_y[177][9] ==1'b1 ? 5'd31 : 
        temp_y[177][3]==1'b1 ? temp_y[177][8:4]+1'b1 : temp_y[177][8:4];
assign temp_y[178] = 
$signed(-{2'b0,x58}<<<3'd1)+$signed({1'b0,x242})+$signed({4'b0,x59}<<<3'd3)+$signed(-{2'b0,x50}<<<3'd1)+$signed(-{2'b0,x251}<<<3'd1)+$signed(-{1'b0,x243})+$signed(-{1'b0,x379})+$signed({1'b0,x114})+$signed(-sharing10)-$signed(11'd8);
assign y178=temp_y[178][11] ==1'b1 ? 5'd0 :  
        temp_y[178][9] ==1'b1 ? 5'd31 : 
        temp_y[178][3]==1'b1 ? temp_y[178][8:4]+1'b1 : temp_y[178][8:4];
assign temp_y[179] = 
$signed(-{1'b0,x122})+$signed({3'b0,x370}<<<3'd2)+$signed(-{2'b0,x50}<<<3'd1)+$signed(-{1'b0,x58})+$signed({3'b0,x378}<<<3'd2)+$signed(-{1'b0,x186})+$signed({2'b0,x179}<<<3'd1)+$signed({2'b0,x59}<<<3'd1)+$signed({1'b0,x187})+$signed(-{2'b0,x250}<<<3'd1)+$signed(-{2'b0,x315}<<<3'd1)+$signed(-{1'b0,x123})+$signed(-{1'b0,x115})+$signed(-{1'b0,x307})+$signed(-{1'b0,x242})+$signed(-{1'b0,x314})+$signed(sharing7)-$signed(11'd16);
assign y179=temp_y[179][11] ==1'b1 ? 5'd0 :  
        temp_y[179][9] ==1'b1 ? 5'd31 : 
        temp_y[179][3]==1'b1 ? temp_y[179][8:4]+1'b1 : temp_y[179][8:4];
assign temp_y[180] = 
$signed(-{1'b0,x369})+$signed(-{4'b0,x314}<<<3'd3)+$signed(-{3'b0,x242}<<<3'd2)+$signed(-{3'b0,x306}<<<3'd2)+$signed(-{1'b0,x377})+$signed(-{4'b0,x307}<<<3'd3)+$signed(-{1'b0,x250})+$signed(-{4'b0,x251}<<<3'd3)+$signed({1'b0,x59})+$signed(-{1'b0,x123})+$signed(-{1'b0,x243})+$signed(-{1'b0,x378})+$signed(-sharing80)+$signed(11'd24);
assign y180=temp_y[180][11] ==1'b1 ? 5'd0 :  
        temp_y[180][9] ==1'b1 ? 5'd31 : 
        temp_y[180][3]==1'b1 ? temp_y[180][8:4]+1'b1 : temp_y[180][8:4];
assign temp_y[181] = 
$signed({1'b0,x114})+$signed({3'b0,x250}<<<3'd2)+$signed({2'b0,x178}<<<3'd1)+$signed({1'b0,x378})+$signed({2'b0,x370}<<<3'd1)+$signed(-{3'b0,x179}<<<3'd2)+$signed(-{2'b0,x314}<<<3'd1)+$signed(-{1'b0,x371})+$signed(-{1'b0,x58})+$signed(-{3'b0,x187}<<<3'd2)+$signed(-{2'b0,x115}<<<3'd1)+$signed(-{1'b0,x307})+$signed({1'b0,x59})+$signed(sharing59)+$signed(11'd16);
assign y181=temp_y[181][11] ==1'b1 ? 5'd0 :  
        temp_y[181][9] ==1'b1 ? 5'd31 : 
        temp_y[181][3]==1'b1 ? temp_y[181][8:4]+1'b1 : temp_y[181][8:4];
assign temp_y[182] = 
$signed(-{1'b0,x125})+$signed(-{3'b0,x380}<<<3'd2)+$signed({2'b0,x316}<<<3'd1)+$signed(-{2'b0,x372}<<<3'd1)+$signed(-{1'b0,x124})+$signed({1'b0,x188})+$signed({2'b0,x309}<<<3'd1)+$signed(-{1'b0,x181})+$signed(-{3'b0,x381}<<<3'd2)+$signed({1'b0,x317})+$signed(sharing41)+$signed(11'd32);
assign y182=temp_y[182][11] ==1'b1 ? 5'd0 :  
        temp_y[182][9] ==1'b1 ? 5'd31 : 
        temp_y[182][3]==1'b1 ? temp_y[182][8:4]+1'b1 : temp_y[182][8:4];
assign temp_y[183] = 
$signed({2'b0,x252}<<<3'd1)+$signed({2'b0,x124}<<<3'd1)+$signed({2'b0,x380}<<<3'd1)+$signed({1'b0,x52})+$signed({1'b0,x116})+$signed(-{1'b0,x309})+$signed(-{1'b0,x316})+$signed(-{2'b0,x253}<<<3'd1)+$signed(-{1'b0,x53})+$signed(-{1'b0,x188})+$signed({3'b0,x381}<<<3'd2)+$signed(sharing41)-$signed(11'd0);
assign y183=temp_y[183][11] ==1'b1 ? 5'd0 :  
        temp_y[183][9] ==1'b1 ? 5'd31 : 
        temp_y[183][3]==1'b1 ? temp_y[183][8:4]+1'b1 : temp_y[183][8:4];
assign temp_y[184] = 
$signed(-{1'b0,x189})+$signed(-{3'b0,x380}<<<3'd2)+$signed(-{2'b0,x372}<<<3'd1)+$signed({2'b0,x252}<<<3'd1)+$signed(-{3'b0,x308}<<<3'd2)+$signed({1'b0,x180})+$signed({1'b0,x244})+$signed(-{2'b0,x116}<<<3'd1)+$signed(-{2'b0,x124}<<<3'd1)+$signed(-{4'b0,x309}<<<3'd3)+$signed(-{3'b0,x316}<<<3'd2)+$signed(-{3'b0,x317}<<<3'd2)+$signed(-{1'b0,x253})+$signed(11'd40);
assign y184=temp_y[184][11] ==1'b1 ? 5'd0 :  
        temp_y[184][9] ==1'b1 ? 5'd31 : 
        temp_y[184][3]==1'b1 ? temp_y[184][8:4]+1'b1 : temp_y[184][8:4];
assign temp_y[185] = 
$signed({2'b0,x372}<<<3'd1)+$signed({1'b0,x308})+$signed({1'b0,x188})+$signed(-{1'b0,x124})+$signed({1'b0,x60})+$signed({1'b0,x373})+$signed(-{2'b0,x125}<<<3'd1)+$signed(-{1'b0,x116})+$signed(-{1'b0,x244})+$signed({1'b0,x317})+$signed(sharing89)+$signed(sharing90)-$signed(11'd16);
assign y185=temp_y[185][11] ==1'b1 ? 5'd0 :  
        temp_y[185][9] ==1'b1 ? 5'd31 : 
        temp_y[185][3]==1'b1 ? temp_y[185][8:4]+1'b1 : temp_y[185][8:4];
assign temp_y[186] = 
$signed({3'b0,x188}<<<3'd2)+$signed(-{2'b0,x60}<<<3'd1)+$signed(-{2'b0,x180}<<<3'd1)+$signed({1'b0,x372})+$signed(-{1'b0,x252})+$signed(-{2'b0,x253}<<<3'd1)+$signed(-{2'b0,x117}<<<3'd1)+$signed(-{2'b0,x373}<<<3'd1)+$signed(sharing89)+$signed(-sharing90)-$signed(11'd24);
assign y186=temp_y[186][11] ==1'b1 ? 5'd0 :  
        temp_y[186][9] ==1'b1 ? 5'd31 : 
        temp_y[186][3]==1'b1 ? temp_y[186][8:4]+1'b1 : temp_y[186][8:4];
assign temp_y[187] = 
$signed(-{1'b0,x381})+$signed({2'b0,x316}<<<3'd1)+$signed({1'b0,x252})+$signed(-{1'b0,x52})+$signed({3'b0,x317}<<<3'd2)+$signed(-{1'b0,x372})+$signed(-{1'b0,x245})+$signed(-{1'b0,x124})+$signed(-{1'b0,x244})+$signed(-{1'b0,x53})+$signed(-sharing26)-$signed(11'd32);
assign y187=temp_y[187][11] ==1'b1 ? 5'd0 :  
        temp_y[187][9] ==1'b1 ? 5'd31 : 
        temp_y[187][3]==1'b1 ? temp_y[187][8:4]+1'b1 : temp_y[187][8:4];
assign temp_y[188] = 
$signed(-{1'b0,x116})+$signed({3'b0,x373}<<<3'd2)+$signed(-{2'b0,x317}<<<3'd1)+$signed({3'b0,x381}<<<3'd2)+$signed(-{2'b0,x309}<<<3'd1)+$signed(-{1'b0,x53})+$signed(-{1'b0,x61})+$signed(sharing64)-$signed(11'd0);
assign y188=temp_y[188][11] ==1'b1 ? 5'd0 :  
        temp_y[188][9] ==1'b1 ? 5'd31 : 
        temp_y[188][3]==1'b1 ? temp_y[188][8:4]+1'b1 : temp_y[188][8:4];
assign temp_y[189] = 
$signed(-{2'b0,x308}<<<3'd1)+$signed({1'b0,x244})+$signed(-{1'b0,x180})+$signed({3'b0,x125}<<<3'd2)+$signed({2'b0,x373}<<<3'd1)+$signed({1'b0,x309})+$signed(-{3'b0,x381}<<<3'd2)+$signed(-{1'b0,x245})+$signed(-{1'b0,x380})+$signed(-sharing112)-$signed(11'd0);
assign y189=temp_y[189][11] ==1'b1 ? 5'd0 :  
        temp_y[189][9] ==1'b1 ? 5'd31 : 
        temp_y[189][3]==1'b1 ? temp_y[189][8:4]+1'b1 : temp_y[189][8:4];
assign temp_y[190] = 
$signed(-{3'b0,x60}<<<3'd2)+$signed(-{2'b0,x244}<<<3'd1)+$signed({1'b0,x380})+$signed(-{1'b0,x316})+$signed(-{1'b0,x188})+$signed({2'b0,x245}<<<3'd1)+$signed(-{2'b0,x61}<<<3'd1)+$signed(-{2'b0,x189}<<<3'd1)+$signed(-{2'b0,x52}<<<3'd1)+$signed({1'b0,x116})+$signed(sharing30)+$signed(11'd40);
assign y190=temp_y[190][11] ==1'b1 ? 5'd0 :  
        temp_y[190][9] ==1'b1 ? 5'd31 : 
        temp_y[190][3]==1'b1 ? temp_y[190][8:4]+1'b1 : temp_y[190][8:4];
assign temp_y[191] = 
$signed(-{2'b0,x60}<<<3'd1)+$signed({1'b0,x244})+$signed({4'b0,x61}<<<3'd3)+$signed(-{1'b0,x245})+$signed(-{2'b0,x253}<<<3'd1)+$signed(-{1'b0,x381})+$signed(-{2'b0,x52}<<<3'd1)+$signed({1'b0,x116})+$signed(-sharing30)-$signed(11'd8);
assign y191=temp_y[191][11] ==1'b1 ? 5'd0 :  
        temp_y[191][9] ==1'b1 ? 5'd31 : 
        temp_y[191][3]==1'b1 ? temp_y[191][8:4]+1'b1 : temp_y[191][8:4];
assign temp_y[192] = 
$signed(-{1'b0,x117})+$signed(-{1'b0,x125})+$signed({1'b0,x189})+$signed({3'b0,x372}<<<3'd2)+$signed({3'b0,x380}<<<3'd2)+$signed(-{2'b0,x52}<<<3'd1)+$signed(-{1'b0,x60})+$signed(-{1'b0,x188})+$signed({2'b0,x181}<<<3'd1)+$signed(-{1'b0,x309})+$signed({2'b0,x61}<<<3'd1)+$signed(-{2'b0,x252}<<<3'd1)+$signed(-{1'b0,x316})+$signed(-{2'b0,x317}<<<3'd1)+$signed(-{1'b0,x124})+$signed(-{1'b0,x244})+$signed(sharing26)-$signed(11'd16);
assign y192=temp_y[192][11] ==1'b1 ? 5'd0 :  
        temp_y[192][9] ==1'b1 ? 5'd31 : 
        temp_y[192][3]==1'b1 ? temp_y[192][8:4]+1'b1 : temp_y[192][8:4];
assign temp_y[193] = 
$signed(-{1'b0,x371})+$signed(-{1'b0,x379})+$signed(-{3'b0,x244}<<<3'd2)+$signed(-{3'b0,x308}<<<3'd2)+$signed(-{4'b0,x316}<<<3'd3)+$signed(-{4'b0,x309}<<<3'd3)+$signed(-{1'b0,x252})+$signed(-{4'b0,x253}<<<3'd3)+$signed(-{1'b0,x125})+$signed(-{1'b0,x245})+$signed(-{1'b0,x380})+$signed({1'b0,x61})+$signed(sharing112)+$signed(11'd24);
assign y193=temp_y[193][11] ==1'b1 ? 5'd0 :  
        temp_y[193][9] ==1'b1 ? 5'd31 : 
        temp_y[193][3]==1'b1 ? temp_y[193][8:4]+1'b1 : temp_y[193][8:4];
assign temp_y[194] = 
$signed(-{1'b0,x309})+$signed({3'b0,x252}<<<3'd2)+$signed({2'b0,x180}<<<3'd1)+$signed({1'b0,x380})+$signed({2'b0,x372}<<<3'd1)+$signed(-{2'b0,x316}<<<3'd1)+$signed(-{1'b0,x60})+$signed(-{1'b0,x373})+$signed(-{3'b0,x181}<<<3'd2)+$signed(-{2'b0,x117}<<<3'd1)+$signed(-{3'b0,x189}<<<3'd2)+$signed({1'b0,x61})+$signed({1'b0,x116})+$signed(sharing64)+$signed(11'd16);
assign y194=temp_y[194][11] ==1'b1 ? 5'd0 :  
        temp_y[194][9] ==1'b1 ? 5'd31 : 
        temp_y[194][3]==1'b1 ? temp_y[194][8:4]+1'b1 : temp_y[194][8:4];
assign temp_y[195] = 
$signed({1'b0,x319})+$signed({2'b0,x318}<<<3'd1)+$signed(-{1'b0,x127})+$signed(-{3'b0,x382}<<<3'd2)+$signed(-{2'b0,x374}<<<3'd1)+$signed(-{1'b0,x126})+$signed({1'b0,x190})+$signed(-{3'b0,x383}<<<3'd2)+$signed({2'b0,x311}<<<3'd1)+$signed(-{1'b0,x183})+$signed(sharing34)+$signed(11'd32);
assign y195=temp_y[195][11] ==1'b1 ? 5'd0 :  
        temp_y[195][9] ==1'b1 ? 5'd31 : 
        temp_y[195][3]==1'b1 ? temp_y[195][8:4]+1'b1 : temp_y[195][8:4];
assign temp_y[196] = 
$signed({2'b0,x254}<<<3'd1)+$signed(-{1'b0,x311})+$signed(-{1'b0,x318})+$signed({2'b0,x382}<<<3'd1)+$signed({1'b0,x118})+$signed({2'b0,x126}<<<3'd1)+$signed({1'b0,x54})+$signed(-{1'b0,x190})+$signed({3'b0,x383}<<<3'd2)+$signed(-{2'b0,x255}<<<3'd1)+$signed(-{1'b0,x55})+$signed(sharing34)-$signed(11'd0);
assign y196=temp_y[196][11] ==1'b1 ? 5'd0 :  
        temp_y[196][9] ==1'b1 ? 5'd31 : 
        temp_y[196][3]==1'b1 ? temp_y[196][8:4]+1'b1 : temp_y[196][8:4];
assign temp_y[197] = 
$signed({2'b0,x254}<<<3'd1)+$signed(-{3'b0,x318}<<<3'd2)+$signed(-{3'b0,x382}<<<3'd2)+$signed(-{2'b0,x118}<<<3'd1)+$signed(-{2'b0,x126}<<<3'd1)+$signed(-{1'b0,x191})+$signed(-{3'b0,x310}<<<3'd2)+$signed(-{2'b0,x374}<<<3'd1)+$signed({1'b0,x246})+$signed(-{4'b0,x311}<<<3'd3)+$signed(-{3'b0,x319}<<<3'd2)+$signed({1'b0,x182})+$signed(-{1'b0,x255})+$signed(11'd40);
assign y197=temp_y[197][11] ==1'b1 ? 5'd0 :  
        temp_y[197][9] ==1'b1 ? 5'd31 : 
        temp_y[197][3]==1'b1 ? temp_y[197][8:4]+1'b1 : temp_y[197][8:4];
assign temp_y[198] = 
$signed({1'b0,x375})+$signed({1'b0,x310})+$signed({1'b0,x62})+$signed(-{1'b0,x118})+$signed(-{1'b0,x126})+$signed({2'b0,x374}<<<3'd1)+$signed(-{1'b0,x246})+$signed({1'b0,x190})+$signed(-{2'b0,x127}<<<3'd1)+$signed({1'b0,x319})+$signed(sharing106)+$signed(sharing107)-$signed(11'd16);
assign y198=temp_y[198][11] ==1'b1 ? 5'd0 :  
        temp_y[198][9] ==1'b1 ? 5'd31 : 
        temp_y[198][3]==1'b1 ? temp_y[198][8:4]+1'b1 : temp_y[198][8:4];
assign temp_y[199] = 
$signed(-{2'b0,x375}<<<3'd1)+$signed(-{2'b0,x62}<<<3'd1)+$signed(-{2'b0,x255}<<<3'd1)+$signed({1'b0,x374})+$signed({3'b0,x190}<<<3'd2)+$signed(-{2'b0,x182}<<<3'd1)+$signed(-{1'b0,x254})+$signed(-{2'b0,x119}<<<3'd1)+$signed(sharing106)+$signed(-sharing107)-$signed(11'd24);
assign y199=temp_y[199][11] ==1'b1 ? 5'd0 :  
        temp_y[199][9] ==1'b1 ? 5'd31 : 
        temp_y[199][3]==1'b1 ? temp_y[199][8:4]+1'b1 : temp_y[199][8:4];
assign temp_y[200] = 
$signed(-{1'b0,x55})+$signed(-{1'b0,x247})+$signed(-{1'b0,x246})+$signed({1'b0,x254})+$signed(-{1'b0,x54})+$signed(-{1'b0,x126})+$signed({2'b0,x318}<<<3'd1)+$signed(-{1'b0,x374})+$signed({3'b0,x319}<<<3'd2)+$signed(-{1'b0,x383})+$signed(sharing23)-$signed(11'd32);
assign y200=temp_y[200][11] ==1'b1 ? 5'd0 :  
        temp_y[200][9] ==1'b1 ? 5'd31 : 
        temp_y[200][3]==1'b1 ? temp_y[200][8:4]+1'b1 : temp_y[200][8:4];
assign temp_y[201] = 
$signed({3'b0,x375}<<<3'd2)+$signed(-{1'b0,x63})+$signed(-{2'b0,x311}<<<3'd1)+$signed(-{1'b0,x118})+$signed({3'b0,x383}<<<3'd2)+$signed(-{2'b0,x319}<<<3'd1)+$signed(-{1'b0,x55})+$signed(sharing52)-$signed(11'd0);
assign y201=temp_y[201][11] ==1'b1 ? 5'd0 :  
        temp_y[201][9] ==1'b1 ? 5'd31 : 
        temp_y[201][3]==1'b1 ? temp_y[201][8:4]+1'b1 : temp_y[201][8:4];
assign temp_y[202] = 
$signed(-{3'b0,x383}<<<3'd2)+$signed(-{1'b0,x247})+$signed({1'b0,x246})+$signed(-{1'b0,x382})+$signed(-{2'b0,x310}<<<3'd1)+$signed(-{1'b0,x182})+$signed({3'b0,x127}<<<3'd2)+$signed({2'b0,x375}<<<3'd1)+$signed({1'b0,x311})+$signed(sharing105)-$signed(11'd0);
assign y202=temp_y[202][11] ==1'b1 ? 5'd0 :  
        temp_y[202][9] ==1'b1 ? 5'd31 : 
        temp_y[202][3]==1'b1 ? temp_y[202][8:4]+1'b1 : temp_y[202][8:4];
assign temp_y[203] = 
$signed(-{2'b0,x54}<<<3'd1)+$signed({1'b0,x382})+$signed({2'b0,x247}<<<3'd1)+$signed(-{2'b0,x63}<<<3'd1)+$signed({1'b0,x118})+$signed(-{3'b0,x62}<<<3'd2)+$signed(-{2'b0,x246}<<<3'd1)+$signed(-{1'b0,x318})+$signed(-{2'b0,x191}<<<3'd1)+$signed(-{1'b0,x190})+$signed(sharing8)+$signed(11'd40);
assign y203=temp_y[203][11] ==1'b1 ? 5'd0 :  
        temp_y[203][9] ==1'b1 ? 5'd31 : 
        temp_y[203][3]==1'b1 ? temp_y[203][8:4]+1'b1 : temp_y[203][8:4];
assign temp_y[204] = 
$signed(-{2'b0,x54}<<<3'd1)+$signed(-{1'b0,x383})+$signed({1'b0,x118})+$signed(-{2'b0,x62}<<<3'd1)+$signed({1'b0,x246})+$signed({4'b0,x63}<<<3'd3)+$signed(-{2'b0,x255}<<<3'd1)+$signed(-{1'b0,x247})+$signed(-sharing8)-$signed(11'd8);
assign y204=temp_y[204][11] ==1'b1 ? 5'd0 :  
        temp_y[204][9] ==1'b1 ? 5'd31 : 
        temp_y[204][3]==1'b1 ? temp_y[204][8:4]+1'b1 : temp_y[204][8:4];
assign temp_y[205] = 
$signed(-{1'b0,x311})+$signed(-{2'b0,x254}<<<3'd1)+$signed(-{1'b0,x246})+$signed(-{1'b0,x119})+$signed({3'b0,x374}<<<3'd2)+$signed({2'b0,x183}<<<3'd1)+$signed(-{1'b0,x62})+$signed({1'b0,x191})+$signed(-{1'b0,x126})+$signed(-{2'b0,x319}<<<3'd1)+$signed({3'b0,x382}<<<3'd2)+$signed(-{2'b0,x54}<<<3'd1)+$signed(-{1'b0,x318})+$signed(-{1'b0,x190})+$signed({2'b0,x63}<<<3'd1)+$signed(-{1'b0,x127})+$signed(-sharing23)-$signed(11'd16);
assign y205=temp_y[205][11] ==1'b1 ? 5'd0 :  
        temp_y[205][9] ==1'b1 ? 5'd31 : 
        temp_y[205][3]==1'b1 ? temp_y[205][8:4]+1'b1 : temp_y[205][8:4];
assign temp_y[206] = 
$signed(-{1'b0,x373})+$signed({1'b0,x63})+$signed(-{3'b0,x310}<<<3'd2)+$signed(-{4'b0,x255}<<<3'd3)+$signed(-{1'b0,x382})+$signed(-{1'b0,x381})+$signed(-{4'b0,x318}<<<3'd3)+$signed(-{3'b0,x246}<<<3'd2)+$signed(-{1'b0,x247})+$signed(-{1'b0,x254})+$signed(-{4'b0,x311}<<<3'd3)+$signed(-{1'b0,x127})+$signed(-sharing105)+$signed(11'd24);
assign y206=temp_y[206][11] ==1'b1 ? 5'd0 :  
        temp_y[206][9] ==1'b1 ? 5'd31 : 
        temp_y[206][3]==1'b1 ? temp_y[206][8:4]+1'b1 : temp_y[206][8:4];
assign temp_y[207] = 
$signed({1'b0,x63})+$signed(-{3'b0,x183}<<<3'd2)+$signed(-{1'b0,x375})+$signed({2'b0,x374}<<<3'd1)+$signed({2'b0,x182}<<<3'd1)+$signed({1'b0,x118})+$signed({1'b0,x382})+$signed({3'b0,x254}<<<3'd2)+$signed(-{2'b0,x318}<<<3'd1)+$signed(-{1'b0,x62})+$signed(-{3'b0,x191}<<<3'd2)+$signed(-{2'b0,x119}<<<3'd1)+$signed(-{1'b0,x311})+$signed(sharing52)+$signed(11'd16);
assign y207=temp_y[207][11] ==1'b1 ? 5'd0 :  
        temp_y[207][9] ==1'b1 ? 5'd31 : 
        temp_y[207][3]==1'b1 ? temp_y[207][8:4]+1'b1 : temp_y[207][8:4];
endmodule