module Conv11(
input [6:0] x0 ,
input [6:0] x1 ,
input [6:0] x2 ,
input [6:0] x3 ,
input [6:0] x4 ,
input [6:0] x5 ,
input [6:0] x6 ,
input [6:0] x7 ,
input [6:0] x8 ,
input [6:0] x9 ,
input [6:0] x10 ,
input [6:0] x11 ,
input [6:0] x12 ,
input [6:0] x13 ,
input [6:0] x14 ,
input [6:0] x15 ,
input [6:0] x16 ,
input [6:0] x17 ,
input [6:0] x18 ,
input [6:0] x19 ,
input [6:0] x20 ,
input [6:0] x21 ,
input [6:0] x22 ,
input [6:0] x23 ,
input [6:0] x24 ,
input [6:0] x25 ,
input [6:0] x26 ,
input [6:0] x27 ,
input [6:0] x28 ,
input [6:0] x29 ,
input [6:0] x30 ,
input [6:0] x31 ,
input [6:0] x32 ,
input [6:0] x33 ,
input [6:0] x34 ,
input [6:0] x35 ,
input [6:0] x36 ,
input [6:0] x37 ,
input [6:0] x38 ,
input [6:0] x39 ,
input [6:0] x40 ,
input [6:0] x41 ,
input [6:0] x42 ,
input [6:0] x43 ,
input [6:0] x44 ,
input [6:0] x45 ,
input [6:0] x46 ,
input [6:0] x47 ,
input [6:0] x48 ,
input [6:0] x49 ,
input [6:0] x50 ,
input [6:0] x51 ,
input [6:0] x52 ,
input [6:0] x53 ,
input [6:0] x54 ,
input [6:0] x55 ,
input [6:0] x56 ,
input [6:0] x57 ,
input [6:0] x58 ,
input [6:0] x59 ,
input [6:0] x60 ,
input [6:0] x61 ,
input [6:0] x62 ,
input [6:0] x63 ,
input [6:0] x64 ,
input [6:0] x65 ,
input [6:0] x66 ,
input [6:0] x67 ,
input [6:0] x68 ,
input [6:0] x69 ,
input [6:0] x70 ,
input [6:0] x71 ,
input [6:0] x72 ,
input [6:0] x73 ,
input [6:0] x74 ,
input [6:0] x75 ,
input [6:0] x76 ,
input [6:0] x77 ,
input [6:0] x78 ,
input [6:0] x79 ,
input [6:0] x80 ,
input [6:0] x81 ,
input [6:0] x82 ,
input [6:0] x83 ,
input [6:0] x84 ,
input [6:0] x85 ,
input [6:0] x86 ,
input [6:0] x87 ,
input [6:0] x88 ,
input [6:0] x89 ,
input [6:0] x90 ,
input [6:0] x91 ,
input [6:0] x92 ,
input [6:0] x93 ,
input [6:0] x94 ,
input [6:0] x95 ,
input [6:0] x96 ,
input [6:0] x97 ,
input [6:0] x98 ,
input [6:0] x99 ,
input [6:0] x100 ,
input [6:0] x101 ,
input [6:0] x102 ,
input [6:0] x103 ,
input [6:0] x104 ,
input [6:0] x105 ,
input [6:0] x106 ,
input [6:0] x107 ,
input [6:0] x108 ,
input [6:0] x109 ,
input [6:0] x110 ,
input [6:0] x111 ,
input [6:0] x112 ,
input [6:0] x113 ,
input [6:0] x114 ,
input [6:0] x115 ,
input [6:0] x116 ,
input [6:0] x117 ,
input [6:0] x118 ,
input [6:0] x119 ,
input [6:0] x120 ,
input [6:0] x121 ,
input [6:0] x122 ,
input [6:0] x123 ,
input [6:0] x124 ,
input [6:0] x125 ,
input [6:0] x126 ,
input [6:0] x127 ,
input [6:0] x128 ,
input [6:0] x129 ,
input [6:0] x130 ,
input [6:0] x131 ,
input [6:0] x132 ,
input [6:0] x133 ,
input [6:0] x134 ,
input [6:0] x135 ,
input [6:0] x136 ,
input [6:0] x137 ,
input [6:0] x138 ,
input [6:0] x139 ,
input [6:0] x140 ,
input [6:0] x141 ,
input [6:0] x142 ,
input [6:0] x143 ,
input [6:0] x144 ,
input [6:0] x145 ,
input [6:0] x146 ,
input [6:0] x147 ,
input [6:0] x148 ,
input [6:0] x149 ,
input [6:0] x150 ,
input [6:0] x151 ,
input [6:0] x152 ,
input [6:0] x153 ,
input [6:0] x154 ,
input [6:0] x155 ,
input [6:0] x156 ,
input [6:0] x157 ,
input [6:0] x158 ,
input [6:0] x159 ,
input [6:0] x160 ,
input [6:0] x161 ,
input [6:0] x162 ,
input [6:0] x163 ,
input [6:0] x164 ,
input [6:0] x165 ,
input [6:0] x166 ,
input [6:0] x167 ,
input [6:0] x168 ,
input [6:0] x169 ,
input [6:0] x170 ,
input [6:0] x171 ,
input [6:0] x172 ,
input [6:0] x173 ,
input [6:0] x174 ,
input [6:0] x175 ,
input [6:0] x176 ,
input [6:0] x177 ,
input [6:0] x178 ,
input [6:0] x179 ,
input [6:0] x180 ,
input [6:0] x181 ,
input [6:0] x182 ,
input [6:0] x183 ,
input [6:0] x184 ,
input [6:0] x185 ,
input [6:0] x186 ,
input [6:0] x187 ,
input [6:0] x188 ,
input [6:0] x189 ,
input [6:0] x190 ,
input [6:0] x191 ,
input [6:0] x192 ,
input [6:0] x193 ,
input [6:0] x194 ,
input [6:0] x195 ,
input [6:0] x196 ,
input [6:0] x197 ,
input [6:0] x198 ,
input [6:0] x199 ,
input [6:0] x200 ,
input [6:0] x201 ,
input [6:0] x202 ,
input [6:0] x203 ,
input [6:0] x204 ,
input [6:0] x205 ,
input [6:0] x206 ,
input [6:0] x207 ,
input [6:0] x208 ,
input [6:0] x209 ,
input [6:0] x210 ,
input [6:0] x211 ,
input [6:0] x212 ,
input [6:0] x213 ,
input [6:0] x214 ,
input [6:0] x215 ,
input [6:0] x216 ,
input [6:0] x217 ,
input [6:0] x218 ,
input [6:0] x219 ,
input [6:0] x220 ,
input [6:0] x221 ,
input [6:0] x222 ,
input [6:0] x223 ,
input [6:0] x224 ,
input [6:0] x225 ,
input [6:0] x226 ,
input [6:0] x227 ,
input [6:0] x228 ,
input [6:0] x229 ,
input [6:0] x230 ,
input [6:0] x231 ,
input [6:0] x232 ,
input [6:0] x233 ,
input [6:0] x234 ,
input [6:0] x235 ,
input [6:0] x236 ,
input [6:0] x237 ,
input [6:0] x238 ,
input [6:0] x239 ,
input [6:0] x240 ,
input [6:0] x241 ,
input [6:0] x242 ,
input [6:0] x243 ,
input [6:0] x244 ,
input [6:0] x245 ,
input [6:0] x246 ,
input [6:0] x247 ,
input [6:0] x248 ,
input [6:0] x249 ,
input [6:0] x250 ,
input [6:0] x251 ,
input [6:0] x252 ,
input [6:0] x253 ,
input [6:0] x254 ,
input [6:0] x255 ,
input [6:0] x256 ,
input [6:0] x257 ,
input [6:0] x258 ,
input [6:0] x259 ,
input [6:0] x260 ,
input [6:0] x261 ,
input [6:0] x262 ,
input [6:0] x263 ,
input [6:0] x264 ,
input [6:0] x265 ,
input [6:0] x266 ,
input [6:0] x267 ,
input [6:0] x268 ,
input [6:0] x269 ,
input [6:0] x270 ,
input [6:0] x271 ,
input [6:0] x272 ,
input [6:0] x273 ,
input [6:0] x274 ,
input [6:0] x275 ,
input [6:0] x276 ,
input [6:0] x277 ,
input [6:0] x278 ,
input [6:0] x279 ,
input [6:0] x280 ,
input [6:0] x281 ,
input [6:0] x282 ,
input [6:0] x283 ,
input [6:0] x284 ,
input [6:0] x285 ,
input [6:0] x286 ,
input [6:0] x287 ,
input [6:0] x288 ,
input [6:0] x289 ,
input [6:0] x290 ,
input [6:0] x291 ,
input [6:0] x292 ,
input [6:0] x293 ,
input [6:0] x294 ,
input [6:0] x295 ,
input [6:0] x296 ,
input [6:0] x297 ,
input [6:0] x298 ,
input [6:0] x299 ,
input [6:0] x300 ,
input [6:0] x301 ,
input [6:0] x302 ,
input [6:0] x303 ,
input [6:0] x304 ,
input [6:0] x305 ,
input [6:0] x306 ,
input [6:0] x307 ,
input [6:0] x308 ,
input [6:0] x309 ,
input [6:0] x310 ,
input [6:0] x311 ,
input [6:0] x312 ,
input [6:0] x313 ,
input [6:0] x314 ,
input [6:0] x315 ,
input [6:0] x316 ,
input [6:0] x317 ,
input [6:0] x318 ,
input [6:0] x319 ,
input [6:0] x320 ,
input [6:0] x321 ,
input [6:0] x322 ,
input [6:0] x323 ,
input [6:0] x324 ,
input [6:0] x325 ,
input [6:0] x326 ,
input [6:0] x327 ,
input [6:0] x328 ,
input [6:0] x329 ,
input [6:0] x330 ,
input [6:0] x331 ,
input [6:0] x332 ,
input [6:0] x333 ,
input [6:0] x334 ,
input [6:0] x335 ,
input [6:0] x336 ,
input [6:0] x337 ,
input [6:0] x338 ,
input [6:0] x339 ,
input [6:0] x340 ,
input [6:0] x341 ,
input [6:0] x342 ,
input [6:0] x343 ,
input [6:0] x344 ,
input [6:0] x345 ,
input [6:0] x346 ,
input [6:0] x347 ,
input [6:0] x348 ,
input [6:0] x349 ,
input [6:0] x350 ,
input [6:0] x351 ,
input [6:0] x352 ,
input [6:0] x353 ,
input [6:0] x354 ,
input [6:0] x355 ,
input [6:0] x356 ,
input [6:0] x357 ,
input [6:0] x358 ,
input [6:0] x359 ,
input [6:0] x360 ,
input [6:0] x361 ,
input [6:0] x362 ,
input [6:0] x363 ,
input [6:0] x364 ,
input [6:0] x365 ,
input [6:0] x366 ,
input [6:0] x367 ,
input [6:0] x368 ,
input [6:0] x369 ,
input [6:0] x370 ,
input [6:0] x371 ,
input [6:0] x372 ,
input [6:0] x373 ,
input [6:0] x374 ,
input [6:0] x375 ,
input [6:0] x376 ,
input [6:0] x377 ,
input [6:0] x378 ,
input [6:0] x379 ,
input [6:0] x380 ,
input [6:0] x381 ,
input [6:0] x382 ,
input [6:0] x383 ,
input [6:0] x384 ,
input [6:0] x385 ,
input [6:0] x386 ,
input [6:0] x387 ,
input [6:0] x388 ,
input [6:0] x389 ,
input [6:0] x390 ,
input [6:0] x391 ,
input [6:0] x392 ,
input [6:0] x393 ,
input [6:0] x394 ,
input [6:0] x395 ,
input [6:0] x396 ,
input [6:0] x397 ,
input [6:0] x398 ,
input [6:0] x399 ,
input [6:0] x400 ,
input [6:0] x401 ,
input [6:0] x402 ,
input [6:0] x403 ,
input [6:0] x404 ,
input [6:0] x405 ,
input [6:0] x406 ,
input [6:0] x407 ,
input [6:0] x408 ,
input [6:0] x409 ,
input [6:0] x410 ,
input [6:0] x411 ,
input [6:0] x412 ,
input [6:0] x413 ,
input [6:0] x414 ,
input [6:0] x415 ,
input [6:0] x416 ,
input [6:0] x417 ,
input [6:0] x418 ,
input [6:0] x419 ,
input [6:0] x420 ,
input [6:0] x421 ,
input [6:0] x422 ,
input [6:0] x423 ,
input [6:0] x424 ,
input [6:0] x425 ,
input [6:0] x426 ,
input [6:0] x427 ,
input [6:0] x428 ,
input [6:0] x429 ,
input [6:0] x430 ,
input [6:0] x431 ,
input [6:0] x432 ,
input [6:0] x433 ,
input [6:0] x434 ,
input [6:0] x435 ,
input [6:0] x436 ,
input [6:0] x437 ,
input [6:0] x438 ,
input [6:0] x439 ,
input [6:0] x440 ,
input [6:0] x441 ,
input [6:0] x442 ,
input [6:0] x443 ,
input [6:0] x444 ,
input [6:0] x445 ,
input [6:0] x446 ,
input [6:0] x447 ,
input [6:0] x448 ,
input [6:0] x449 ,
input [6:0] x450 ,
input [6:0] x451 ,
input [6:0] x452 ,
input [6:0] x453 ,
input [6:0] x454 ,
input [6:0] x455 ,
input [6:0] x456 ,
input [6:0] x457 ,
input [6:0] x458 ,
input [6:0] x459 ,
input [6:0] x460 ,
input [6:0] x461 ,
input [6:0] x462 ,
input [6:0] x463 ,
input [6:0] x464 ,
input [6:0] x465 ,
input [6:0] x466 ,
input [6:0] x467 ,
input [6:0] x468 ,
input [6:0] x469 ,
input [6:0] x470 ,
input [6:0] x471 ,
input [6:0] x472 ,
input [6:0] x473 ,
input [6:0] x474 ,
input [6:0] x475 ,
input [6:0] x476 ,
input [6:0] x477 ,
input [6:0] x478 ,
input [6:0] x479 ,
input [6:0] x480 ,
input [6:0] x481 ,
input [6:0] x482 ,
input [6:0] x483 ,
input [6:0] x484 ,
input [6:0] x485 ,
input [6:0] x486 ,
input [6:0] x487 ,
input [6:0] x488 ,
input [6:0] x489 ,
input [6:0] x490 ,
input [6:0] x491 ,
input [6:0] x492 ,
input [6:0] x493 ,
input [6:0] x494 ,
input [6:0] x495 ,
input [6:0] x496 ,
input [6:0] x497 ,
input [6:0] x498 ,
input [6:0] x499 ,
input [6:0] x500 ,
input [6:0] x501 ,
input [6:0] x502 ,
input [6:0] x503 ,
input [6:0] x504 ,
input [6:0] x505 ,
input [6:0] x506 ,
input [6:0] x507 ,
input [6:0] x508 ,
input [6:0] x509 ,
input [6:0] x510 ,
input [6:0] x511 ,
input [6:0] x512 ,
input [6:0] x513 ,
input [6:0] x514 ,
input [6:0] x515 ,
input [6:0] x516 ,
input [6:0] x517 ,
input [6:0] x518 ,
input [6:0] x519 ,
input [6:0] x520 ,
input [6:0] x521 ,
input [6:0] x522 ,
input [6:0] x523 ,
input [6:0] x524 ,
input [6:0] x525 ,
input [6:0] x526 ,
input [6:0] x527 ,
input [6:0] x528 ,
input [6:0] x529 ,
input [6:0] x530 ,
input [6:0] x531 ,
input [6:0] x532 ,
input [6:0] x533 ,
input [6:0] x534 ,
input [6:0] x535 ,
input [6:0] x536 ,
input [6:0] x537 ,
input [6:0] x538 ,
input [6:0] x539 ,
input [6:0] x540 ,
input [6:0] x541 ,
input [6:0] x542 ,
input [6:0] x543 ,
input [6:0] x544 ,
input [6:0] x545 ,
input [6:0] x546 ,
input [6:0] x547 ,
input [6:0] x548 ,
input [6:0] x549 ,
input [6:0] x550 ,
input [6:0] x551 ,
input [6:0] x552 ,
input [6:0] x553 ,
input [6:0] x554 ,
input [6:0] x555 ,
input [6:0] x556 ,
input [6:0] x557 ,
input [6:0] x558 ,
input [6:0] x559 ,
input [6:0] x560 ,
input [6:0] x561 ,
input [6:0] x562 ,
input [6:0] x563 ,
input [6:0] x564 ,
input [6:0] x565 ,
input [6:0] x566 ,
input [6:0] x567 ,
input [6:0] x568 ,
input [6:0] x569 ,
input [6:0] x570 ,
input [6:0] x571 ,
input [6:0] x572 ,
input [6:0] x573 ,
input [6:0] x574 ,
input [6:0] x575 ,
input [6:0] x576 ,
input [6:0] x577 ,
input [6:0] x578 ,
input [6:0] x579 ,
input [6:0] x580 ,
input [6:0] x581 ,
input [6:0] x582 ,
input [6:0] x583 ,
input [6:0] x584 ,
input [6:0] x585 ,
input [6:0] x586 ,
input [6:0] x587 ,
input [6:0] x588 ,
input [6:0] x589 ,
input [6:0] x590 ,
input [6:0] x591 ,
input [6:0] x592 ,
input [6:0] x593 ,
input [6:0] x594 ,
input [6:0] x595 ,
input [6:0] x596 ,
input [6:0] x597 ,
input [6:0] x598 ,
input [6:0] x599 ,
input [6:0] x600 ,
input [6:0] x601 ,
input [6:0] x602 ,
input [6:0] x603 ,
input [6:0] x604 ,
input [6:0] x605 ,
input [6:0] x606 ,
input [6:0] x607 ,
input [6:0] x608 ,
input [6:0] x609 ,
input [6:0] x610 ,
input [6:0] x611 ,
input [6:0] x612 ,
input [6:0] x613 ,
input [6:0] x614 ,
input [6:0] x615 ,
input [6:0] x616 ,
input [6:0] x617 ,
input [6:0] x618 ,
input [6:0] x619 ,
input [6:0] x620 ,
input [6:0] x621 ,
input [6:0] x622 ,
input [6:0] x623 ,
input [6:0] x624 ,
input [6:0] x625 ,
input [6:0] x626 ,
input [6:0] x627 ,
input [6:0] x628 ,
input [6:0] x629 ,
input [6:0] x630 ,
input [6:0] x631 ,
input [6:0] x632 ,
input [6:0] x633 ,
input [6:0] x634 ,
input [6:0] x635 ,
input [6:0] x636 ,
input [6:0] x637 ,
input [6:0] x638 ,
input [6:0] x639 ,
input [6:0] x640 ,
input [6:0] x641 ,
input [6:0] x642 ,
input [6:0] x643 ,
input [6:0] x644 ,
input [6:0] x645 ,
input [6:0] x646 ,
input [6:0] x647 ,
input [6:0] x648 ,
input [6:0] x649 ,
input [6:0] x650 ,
input [6:0] x651 ,
input [6:0] x652 ,
input [6:0] x653 ,
input [6:0] x654 ,
input [6:0] x655 ,
input [6:0] x656 ,
input [6:0] x657 ,
input [6:0] x658 ,
input [6:0] x659 ,
input [6:0] x660 ,
input [6:0] x661 ,
input [6:0] x662 ,
input [6:0] x663 ,
input [6:0] x664 ,
input [6:0] x665 ,
input [6:0] x666 ,
input [6:0] x667 ,
input [6:0] x668 ,
input [6:0] x669 ,
input [6:0] x670 ,
input [6:0] x671 ,
input [6:0] x672 ,
input [6:0] x673 ,
input [6:0] x674 ,
input [6:0] x675 ,
input [6:0] x676 ,
input [6:0] x677 ,
input [6:0] x678 ,
input [6:0] x679 ,
input [6:0] x680 ,
input [6:0] x681 ,
input [6:0] x682 ,
input [6:0] x683 ,
input [6:0] x684 ,
input [6:0] x685 ,
input [6:0] x686 ,
input [6:0] x687 ,
input [6:0] x688 ,
input [6:0] x689 ,
input [6:0] x690 ,
input [6:0] x691 ,
input [6:0] x692 ,
input [6:0] x693 ,
input [6:0] x694 ,
input [6:0] x695 ,
input [6:0] x696 ,
input [6:0] x697 ,
input [6:0] x698 ,
input [6:0] x699 ,
input [6:0] x700 ,
input [6:0] x701 ,
input [6:0] x702 ,
input [6:0] x703 ,
input [6:0] x704 ,
input [6:0] x705 ,
input [6:0] x706 ,
input [6:0] x707 ,
input [6:0] x708 ,
input [6:0] x709 ,
input [6:0] x710 ,
input [6:0] x711 ,
input [6:0] x712 ,
input [6:0] x713 ,
input [6:0] x714 ,
input [6:0] x715 ,
input [6:0] x716 ,
input [6:0] x717 ,
input [6:0] x718 ,
input [6:0] x719 ,
input [6:0] x720 ,
input [6:0] x721 ,
input [6:0] x722 ,
input [6:0] x723 ,
input [6:0] x724 ,
input [6:0] x725 ,
input [6:0] x726 ,
input [6:0] x727 ,
input [6:0] x728 ,
input [6:0] x729 ,
input [6:0] x730 ,
input [6:0] x731 ,
input [6:0] x732 ,
input [6:0] x733 ,
input [6:0] x734 ,
input [6:0] x735 ,
input [6:0] x736 ,
input [6:0] x737 ,
input [6:0] x738 ,
input [6:0] x739 ,
input [6:0] x740 ,
input [6:0] x741 ,
input [6:0] x742 ,
input [6:0] x743 ,
input [6:0] x744 ,
input [6:0] x745 ,
input [6:0] x746 ,
input [6:0] x747 ,
input [6:0] x748 ,
input [6:0] x749 ,
input [6:0] x750 ,
input [6:0] x751 ,
input [6:0] x752 ,
input [6:0] x753 ,
input [6:0] x754 ,
input [6:0] x755 ,
input [6:0] x756 ,
input [6:0] x757 ,
input [6:0] x758 ,
input [6:0] x759 ,
input [6:0] x760 ,
input [6:0] x761 ,
input [6:0] x762 ,
input [6:0] x763 ,
input [6:0] x764 ,
input [6:0] x765 ,
input [6:0] x766 ,
input [6:0] x767 ,
output [4:0] y0 ,
output [4:0] y1 ,
output [4:0] y2 ,
output [4:0] y3 ,
output [4:0] y4 ,
output [4:0] y5 ,
output [4:0] y6 ,
output [4:0] y7 ,
output [4:0] y8 ,
output [4:0] y9 ,
output [4:0] y10 ,
output [4:0] y11 ,
output [4:0] y12 ,
output [4:0] y13 ,
output [4:0] y14 ,
output [4:0] y15 ,
output [4:0] y16 ,
output [4:0] y17 ,
output [4:0] y18 ,
output [4:0] y19 ,
output [4:0] y20 ,
output [4:0] y21 ,
output [4:0] y22 ,
output [4:0] y23 ,
output [4:0] y24 ,
output [4:0] y25 ,
output [4:0] y26 ,
output [4:0] y27 ,
output [4:0] y28 ,
output [4:0] y29 ,
output [4:0] y30 ,
output [4:0] y31 ,
output [4:0] y32 ,
output [4:0] y33 ,
output [4:0] y34 ,
output [4:0] y35 ,
output [4:0] y36 ,
output [4:0] y37 ,
output [4:0] y38 ,
output [4:0] y39 ,
output [4:0] y40 ,
output [4:0] y41 ,
output [4:0] y42 ,
output [4:0] y43 ,
output [4:0] y44 ,
output [4:0] y45 ,
output [4:0] y46 ,
output [4:0] y47 ,
output [4:0] y48 ,
output [4:0] y49 ,
output [4:0] y50 ,
output [4:0] y51 ,
output [4:0] y52 ,
output [4:0] y53 ,
output [4:0] y54 ,
output [4:0] y55 ,
output [4:0] y56 ,
output [4:0] y57 ,
output [4:0] y58 ,
output [4:0] y59 ,
output [4:0] y60 ,
output [4:0] y61 ,
output [4:0] y62 ,
output [4:0] y63 ,
output [4:0] y64 ,
output [4:0] y65 ,
output [4:0] y66 ,
output [4:0] y67 ,
output [4:0] y68 ,
output [4:0] y69 ,
output [4:0] y70 ,
output [4:0] y71 ,
output [4:0] y72 ,
output [4:0] y73 ,
output [4:0] y74 ,
output [4:0] y75 ,
output [4:0] y76 ,
output [4:0] y77 ,
output [4:0] y78 ,
output [4:0] y79 ,
output [4:0] y80 ,
output [4:0] y81 ,
output [4:0] y82 ,
output [4:0] y83 ,
output [4:0] y84 ,
output [4:0] y85 ,
output [4:0] y86 ,
output [4:0] y87 ,
output [4:0] y88 ,
output [4:0] y89 ,
output [4:0] y90 ,
output [4:0] y91 ,
output [4:0] y92 ,
output [4:0] y93 ,
output [4:0] y94 ,
output [4:0] y95 ,
output [4:0] y96 ,
output [4:0] y97 ,
output [4:0] y98 ,
output [4:0] y99 ,
output [4:0] y100 ,
output [4:0] y101 ,
output [4:0] y102 ,
output [4:0] y103 ,
output [4:0] y104 ,
output [4:0] y105 ,
output [4:0] y106 ,
output [4:0] y107 ,
output [4:0] y108 ,
output [4:0] y109 ,
output [4:0] y110 ,
output [4:0] y111 ,
output [4:0] y112 ,
output [4:0] y113 ,
output [4:0] y114 ,
output [4:0] y115 ,
output [4:0] y116 ,
output [4:0] y117 ,
output [4:0] y118 ,
output [4:0] y119 ,
output [4:0] y120 ,
output [4:0] y121 ,
output [4:0] y122 ,
output [4:0] y123 ,
output [4:0] y124 ,
output [4:0] y125 ,
output [4:0] y126 ,
output [4:0] y127 ,
output [4:0] y128 ,
output [4:0] y129 ,
output [4:0] y130 ,
output [4:0] y131 ,
output [4:0] y132 ,
output [4:0] y133 ,
output [4:0] y134 ,
output [4:0] y135 ,
output [4:0] y136 ,
output [4:0] y137 ,
output [4:0] y138 ,
output [4:0] y139 ,
output [4:0] y140 ,
output [4:0] y141 ,
output [4:0] y142 ,
output [4:0] y143 ,
output [4:0] y144 ,
output [4:0] y145 ,
output [4:0] y146 ,
output [4:0] y147 ,
output [4:0] y148 ,
output [4:0] y149 ,
output [4:0] y150 ,
output [4:0] y151 ,
output [4:0] y152 ,
output [4:0] y153 ,
output [4:0] y154 ,
output [4:0] y155 ,
output [4:0] y156 ,
output [4:0] y157 ,
output [4:0] y158 ,
output [4:0] y159 ,
output [4:0] y160 ,
output [4:0] y161 ,
output [4:0] y162 ,
output [4:0] y163 ,
output [4:0] y164 ,
output [4:0] y165 ,
output [4:0] y166 ,
output [4:0] y167 ,
output [4:0] y168 ,
output [4:0] y169 ,
output [4:0] y170 ,
output [4:0] y171 ,
output [4:0] y172 ,
output [4:0] y173 ,
output [4:0] y174 ,
output [4:0] y175 ,
output [4:0] y176 ,
output [4:0] y177 ,
output [4:0] y178 ,
output [4:0] y179 ,
output [4:0] y180 ,
output [4:0] y181 ,
output [4:0] y182 ,
output [4:0] y183 ,
output [4:0] y184 ,
output [4:0] y185 ,
output [4:0] y186 ,
output [4:0] y187 ,
output [4:0] y188 ,
output [4:0] y189 ,
output [4:0] y190 ,
output [4:0] y191 ,
output [4:0] y192 ,
output [4:0] y193 ,
output [4:0] y194 ,
output [4:0] y195 ,
output [4:0] y196 ,
output [4:0] y197 ,
output [4:0] y198 ,
output [4:0] y199 ,
output [4:0] y200 ,
output [4:0] y201 ,
output [4:0] y202 ,
output [4:0] y203 ,
output [4:0] y204 ,
output [4:0] y205 ,
output [4:0] y206 ,
output [4:0] y207 ,
output [4:0] y208 ,
output [4:0] y209 ,
output [4:0] y210 ,
output [4:0] y211 ,
output [4:0] y212 ,
output [4:0] y213 ,
output [4:0] y214 ,
output [4:0] y215 ,
output [4:0] y216 ,
output [4:0] y217 ,
output [4:0] y218 ,
output [4:0] y219 ,
output [4:0] y220 ,
output [4:0] y221 ,
output [4:0] y222 ,
output [4:0] y223 ,
output [4:0] y224 ,
output [4:0] y225 ,
output [4:0] y226 ,
output [4:0] y227 ,
output [4:0] y228 ,
output [4:0] y229 ,
output [4:0] y230 ,
output [4:0] y231 ,
output [4:0] y232 ,
output [4:0] y233 ,
output [4:0] y234 ,
output [4:0] y235 ,
output [4:0] y236 ,
output [4:0] y237 ,
output [4:0] y238 ,
output [4:0] y239 ,
output [4:0] y240 ,
output [4:0] y241 ,
output [4:0] y242 ,
output [4:0] y243 ,
output [4:0] y244 ,
output [4:0] y245 ,
output [4:0] y246 ,
output [4:0] y247 ,
output [4:0] y248 ,
output [4:0] y249 ,
output [4:0] y250 ,
output [4:0] y251 ,
output [4:0] y252 ,
output [4:0] y253 ,
output [4:0] y254 ,
output [4:0] y255 ,
output [4:0] y256 ,
output [4:0] y257 ,
output [4:0] y258 ,
output [4:0] y259 ,
output [4:0] y260 ,
output [4:0] y261 ,
output [4:0] y262 ,
output [4:0] y263 ,
output [4:0] y264 ,
output [4:0] y265 ,
output [4:0] y266 ,
output [4:0] y267 ,
output [4:0] y268 ,
output [4:0] y269 ,
output [4:0] y270 ,
output [4:0] y271 ,
output [4:0] y272 ,
output [4:0] y273 ,
output [4:0] y274 ,
output [4:0] y275 ,
output [4:0] y276 ,
output [4:0] y277 ,
output [4:0] y278 ,
output [4:0] y279 ,
output [4:0] y280 ,
output [4:0] y281 ,
output [4:0] y282 ,
output [4:0] y283 ,
output [4:0] y284 ,
output [4:0] y285 ,
output [4:0] y286 ,
output [4:0] y287 ,
output [4:0] y288 ,
output [4:0] y289 ,
output [4:0] y290 ,
output [4:0] y291 ,
output [4:0] y292 ,
output [4:0] y293 ,
output [4:0] y294 ,
output [4:0] y295 ,
output [4:0] y296 ,
output [4:0] y297 ,
output [4:0] y298 ,
output [4:0] y299 ,
output [4:0] y300 ,
output [4:0] y301 ,
output [4:0] y302 ,
output [4:0] y303 ,
output [4:0] y304 ,
output [4:0] y305 ,
output [4:0] y306 ,
output [4:0] y307 ,
output [4:0] y308 ,
output [4:0] y309 ,
output [4:0] y310 ,
output [4:0] y311 ,
output [4:0] y312 ,
output [4:0] y313 ,
output [4:0] y314 ,
output [4:0] y315 ,
output [4:0] y316 ,
output [4:0] y317 ,
output [4:0] y318 ,
output [4:0] y319 ,
output [4:0] y320 ,
output [4:0] y321 ,
output [4:0] y322 ,
output [4:0] y323 ,
output [4:0] y324 ,
output [4:0] y325 ,
output [4:0] y326 ,
output [4:0] y327 ,
output [4:0] y328 ,
output [4:0] y329 ,
output [4:0] y330 ,
output [4:0] y331 ,
output [4:0] y332 ,
output [4:0] y333 ,
output [4:0] y334 ,
output [4:0] y335 ,
output [4:0] y336 ,
output [4:0] y337 ,
output [4:0] y338 ,
output [4:0] y339 ,
output [4:0] y340 ,
output [4:0] y341 ,
output [4:0] y342 ,
output [4:0] y343 ,
output [4:0] y344 ,
output [4:0] y345 ,
output [4:0] y346 ,
output [4:0] y347 ,
output [4:0] y348 ,
output [4:0] y349 ,
output [4:0] y350 ,
output [4:0] y351 ,
output [4:0] y352 ,
output [4:0] y353 ,
output [4:0] y354 ,
output [4:0] y355 ,
output [4:0] y356 ,
output [4:0] y357 ,
output [4:0] y358 ,
output [4:0] y359 ,
output [4:0] y360 ,
output [4:0] y361 ,
output [4:0] y362 ,
output [4:0] y363 ,
output [4:0] y364 ,
output [4:0] y365 ,
output [4:0] y366 ,
output [4:0] y367 ,
output [4:0] y368 ,
output [4:0] y369 ,
output [4:0] y370 ,
output [4:0] y371 ,
output [4:0] y372 ,
output [4:0] y373 ,
output [4:0] y374 ,
output [4:0] y375 ,
output [4:0] y376 ,
output [4:0] y377 ,
output [4:0] y378 ,
output [4:0] y379 ,
output [4:0] y380 ,
output [4:0] y381 ,
output [4:0] y382 ,
output [4:0] y383 ,
output [4:0] y384 ,
output [4:0] y385 ,
output [4:0] y386 ,
output [4:0] y387 ,
output [4:0] y388 ,
output [4:0] y389 ,
output [4:0] y390 ,
output [4:0] y391 ,
output [4:0] y392 ,
output [4:0] y393 ,
output [4:0] y394 ,
output [4:0] y395 ,
output [4:0] y396 ,
output [4:0] y397 ,
output [4:0] y398 ,
output [4:0] y399 ,
output [4:0] y400 ,
output [4:0] y401 ,
output [4:0] y402 ,
output [4:0] y403 ,
output [4:0] y404 ,
output [4:0] y405 ,
output [4:0] y406 ,
output [4:0] y407 ,
output [4:0] y408 ,
output [4:0] y409 ,
output [4:0] y410 ,
output [4:0] y411 ,
output [4:0] y412 ,
output [4:0] y413 ,
output [4:0] y414 ,
output [4:0] y415 ,
output [4:0] y416 ,
output [4:0] y417 ,
output [4:0] y418 ,
output [4:0] y419 ,
output [4:0] y420 ,
output [4:0] y421 ,
output [4:0] y422 ,
output [4:0] y423 ,
output [4:0] y424 ,
output [4:0] y425 ,
output [4:0] y426 ,
output [4:0] y427 ,
output [4:0] y428 ,
output [4:0] y429 ,
output [4:0] y430 ,
output [4:0] y431 ,
output [4:0] y432 ,
output [4:0] y433 ,
output [4:0] y434 ,
output [4:0] y435 ,
output [4:0] y436 ,
output [4:0] y437 ,
output [4:0] y438 ,
output [4:0] y439 ,
output [4:0] y440 ,
output [4:0] y441 ,
output [4:0] y442 ,
output [4:0] y443 ,
output [4:0] y444 ,
output [4:0] y445 ,
output [4:0] y446 ,
output [4:0] y447 ,
output [4:0] y448 ,
output [4:0] y449 ,
output [4:0] y450 ,
output [4:0] y451 ,
output [4:0] y452 ,
output [4:0] y453 ,
output [4:0] y454 ,
output [4:0] y455 ,
output [4:0] y456 ,
output [4:0] y457 ,
output [4:0] y458 ,
output [4:0] y459 ,
output [4:0] y460 ,
output [4:0] y461 ,
output [4:0] y462 ,
output [4:0] y463 ,
output [4:0] y464 ,
output [4:0] y465 ,
output [4:0] y466 ,
output [4:0] y467 ,
output [4:0] y468 ,
output [4:0] y469 ,
output [4:0] y470 ,
output [4:0] y471 ,
output [4:0] y472 ,
output [4:0] y473 ,
output [4:0] y474 ,
output [4:0] y475 ,
output [4:0] y476 ,
output [4:0] y477 ,
output [4:0] y478 ,
output [4:0] y479 ,
output [4:0] y480 ,
output [4:0] y481 ,
output [4:0] y482 ,
output [4:0] y483 ,
output [4:0] y484 ,
output [4:0] y485 ,
output [4:0] y486 ,
output [4:0] y487 ,
output [4:0] y488 ,
output [4:0] y489 ,
output [4:0] y490 ,
output [4:0] y491 ,
output [4:0] y492 ,
output [4:0] y493 ,
output [4:0] y494 ,
output [4:0] y495 ,
output [4:0] y496 ,
output [4:0] y497 ,
output [4:0] y498 ,
output [4:0] y499 ,
output [4:0] y500 ,
output [4:0] y501 ,
output [4:0] y502 ,
output [4:0] y503 ,
output [4:0] y504 ,
output [4:0] y505 ,
output [4:0] y506 ,
output [4:0] y507 ,
output [4:0] y508 ,
output [4:0] y509 ,
output [4:0] y510 ,
output [4:0] y511 ,
output [4:0] y512 ,
output [4:0] y513 ,
output [4:0] y514 ,
output [4:0] y515 ,
output [4:0] y516 ,
output [4:0] y517 ,
output [4:0] y518 ,
output [4:0] y519 ,
output [4:0] y520 ,
output [4:0] y521 ,
output [4:0] y522 ,
output [4:0] y523 ,
output [4:0] y524 ,
output [4:0] y525 ,
output [4:0] y526 ,
output [4:0] y527 ,
output [4:0] y528 ,
output [4:0] y529 ,
output [4:0] y530 ,
output [4:0] y531 ,
output [4:0] y532 ,
output [4:0] y533 ,
output [4:0] y534 ,
output [4:0] y535 ,
output [4:0] y536 ,
output [4:0] y537 ,
output [4:0] y538 ,
output [4:0] y539 ,
output [4:0] y540 ,
output [4:0] y541 ,
output [4:0] y542 ,
output [4:0] y543 ,
output [4:0] y544 ,
output [4:0] y545 ,
output [4:0] y546 ,
output [4:0] y547 ,
output [4:0] y548 ,
output [4:0] y549 ,
output [4:0] y550 ,
output [4:0] y551 ,
output [4:0] y552 ,
output [4:0] y553 ,
output [4:0] y554 ,
output [4:0] y555 ,
output [4:0] y556 ,
output [4:0] y557 ,
output [4:0] y558 ,
output [4:0] y559 ,
output [4:0] y560 ,
output [4:0] y561 ,
output [4:0] y562 ,
output [4:0] y563 ,
output [4:0] y564 ,
output [4:0] y565 ,
output [4:0] y566 ,
output [4:0] y567 ,
output [4:0] y568 ,
output [4:0] y569 ,
output [4:0] y570 ,
output [4:0] y571 ,
output [4:0] y572 ,
output [4:0] y573 ,
output [4:0] y574 ,
output [4:0] y575 ,
output [4:0] y576 ,
output [4:0] y577 ,
output [4:0] y578 ,
output [4:0] y579 ,
output [4:0] y580 ,
output [4:0] y581 ,
output [4:0] y582 ,
output [4:0] y583 ,
output [4:0] y584 ,
output [4:0] y585 ,
output [4:0] y586 ,
output [4:0] y587 ,
output [4:0] y588 ,
output [4:0] y589 ,
output [4:0] y590 ,
output [4:0] y591 ,
output [4:0] y592 ,
output [4:0] y593 ,
output [4:0] y594 ,
output [4:0] y595 ,
output [4:0] y596 ,
output [4:0] y597 ,
output [4:0] y598 ,
output [4:0] y599 ,
output [4:0] y600 ,
output [4:0] y601 ,
output [4:0] y602 ,
output [4:0] y603 ,
output [4:0] y604 ,
output [4:0] y605 ,
output [4:0] y606 ,
output [4:0] y607 ,
output [4:0] y608 ,
output [4:0] y609 ,
output [4:0] y610 ,
output [4:0] y611 ,
output [4:0] y612 ,
output [4:0] y613 ,
output [4:0] y614 ,
output [4:0] y615 ,
output [4:0] y616 ,
output [4:0] y617 ,
output [4:0] y618 ,
output [4:0] y619 ,
output [4:0] y620 ,
output [4:0] y621 ,
output [4:0] y622 ,
output [4:0] y623 ,
output [4:0] y624 ,
output [4:0] y625 ,
output [4:0] y626 ,
output [4:0] y627 ,
output [4:0] y628 ,
output [4:0] y629 ,
output [4:0] y630 ,
output [4:0] y631 ,
output [4:0] y632 ,
output [4:0] y633 ,
output [4:0] y634 ,
output [4:0] y635 ,
output [4:0] y636 ,
output [4:0] y637 ,
output [4:0] y638 ,
output [4:0] y639 
);
wire signed[11:0] temp_y  [0:639];
assign temp_y[0] = 
+$signed( -{ 2'b0,x256 }<<<3'd1 )+$signed( -{ 1'b0,x512 } )+$signed( { 1'b0,x1 }  )+$signed( { 1'b0,x257 }  )+$signed( { 1'b0,x513 }  )+$signed( -{ 2'b0,x272 }<<<3'd1 )+$signed( -{ 2'b0,x528 }<<<3'd1 )+$signed( { 2'b0,x273 } <<<3'd1 )+$signed( { 2'b0,x529 } <<<3'd1 )-$signed(11'd16);
assign y0=temp_y[0][11] ==1'b1 ? 5'd0 :  
        temp_y[0][8] ==1'b1 ? 5'd31 : 
        temp_y[0][2]==1'b1 ? temp_y[0][7:3]+1'b1 : temp_y[0][7:3];
assign temp_y[64] = 
+$signed( { 3'b0,x0 }<<<3'd2 )+$signed( -{ 2'b0,x256 }<<<3'd1 )+$signed( -{ 2'b0,x512 }<<<3'd1 )+$signed( { 2'b0,x1 } <<<3'd1 )+$signed( -{ 3'b0,x257 }<<<3'd2)+$signed( { 1'b0,x513 }  )+$signed( -{ 1'b0,x16 } )+$signed( { 1'b0,x528 }  )+$signed( -{ 2'b0,x17 }<<<3'd1 )+$signed( -{ 1'b0,x273 } )+$signed( { 2'b0,x529 } <<<3'd1 )+$signed(11'd24);
assign y64=temp_y[64][11] ==1'b1 ? 5'd0 :  
        temp_y[64][8] ==1'b1 ? 5'd31 : 
        temp_y[64][2]==1'b1 ? temp_y[64][7:3]+1'b1 : temp_y[64][7:3];
assign temp_y[128] = 
+$signed( { 2'b0,x0 } <<<3'd1 )+$signed( { 2'b0,x256 } <<<3'd1 )+$signed( { 1'b0,x512 }  )+$signed( { 2'b0,x1 } <<<3'd1 )+$signed( -{ 1'b0,x257 } )+$signed( { 1'b0,x513 }  )+$signed( -{ 2'b0,x16 }<<<3'd1 )+$signed( -{ 2'b0,x272 }<<<3'd1 )+$signed( -{ 1'b0,x528 } )+$signed( -{ 1'b0,x17 } )+$signed( -{ 1'b0,x273 } )+$signed( -{ 1'b0,x529 } )+$signed(11'd16);
assign y128=temp_y[128][11] ==1'b1 ? 5'd0 :  
        temp_y[128][8] ==1'b1 ? 5'd31 : 
        temp_y[128][2]==1'b1 ? temp_y[128][7:3]+1'b1 : temp_y[128][7:3];
assign temp_y[192] = 
+$signed( { 1'b0,x0 }  )+$signed( -{ 1'b0,x256 } )+$signed( { 1'b0,x1 }  )+$signed( -{ 1'b0,x257 } )+$signed( { 2'b0,x16 } <<<3'd1 )+$signed( -{ 1'b0,x272 } )+$signed( -{ 1'b0,x528 } )+$signed( { 2'b0,x17 } <<<3'd1 )+$signed( -{ 1'b0,x273 } )+$signed( -{ 2'b0,x529 }<<<3'd1 )+$signed(11'd40);
assign y192=temp_y[192][11] ==1'b1 ? 5'd0 :  
        temp_y[192][8] ==1'b1 ? 5'd31 : 
        temp_y[192][2]==1'b1 ? temp_y[192][7:3]+1'b1 : temp_y[192][7:3];
assign temp_y[256] = 
+$signed( -{ 1'b0,x0 } )+$signed( { 2'b0,x256 } <<<3'd1 )+$signed( -{ 1'b0,x512 } )+$signed( -{ 1'b0,x1 } )+$signed( { 2'b0,x257 } <<<3'd1 )+$signed( -{ 2'b0,x513 }<<<3'd1 )+$signed( -{ 1'b0,x16 } )+$signed( { 2'b0,x272 } <<<3'd1 )+$signed( -{ 1'b0,x528 } )+$signed( -{ 2'b0,x17 }<<<3'd1 )+$signed( { 3'b0,x273 }<<<3'd2 )+$signed( -{ 2'b0,x529 }<<<3'd1 )+$signed(11'd32);
assign y256=temp_y[256][11] ==1'b1 ? 5'd0 :  
        temp_y[256][8] ==1'b1 ? 5'd31 : 
        temp_y[256][2]==1'b1 ? temp_y[256][7:3]+1'b1 : temp_y[256][7:3];
assign temp_y[320] = 
+$signed( -{ 1'b0,x0 } )+$signed( -{ 2'b0,x256 }<<<3'd1 )+$signed( -{ 1'b0,x512 } )+$signed( { 1'b0,x1 }  )+$signed( { 2'b0,x257 } <<<3'd1 )+$signed( { 1'b0,x513 }  )+$signed( { 1'b0,x16 }  )+$signed( { 2'b0,x272 } <<<3'd1 )+$signed( { 2'b0,x528 } <<<3'd1 )+$signed( -{ 1'b0,x17 } )+$signed( -{ 2'b0,x273 }<<<3'd1 )+$signed( -{ 1'b0,x529 } )-$signed(11'd68);
assign y320=temp_y[320][11] ==1'b1 ? 5'd0 :  
        temp_y[320][8] ==1'b1 ? 5'd31 : 
        temp_y[320][2]==1'b1 ? temp_y[320][7:3]+1'b1 : temp_y[320][7:3];
assign temp_y[384] = 
+$signed( { 1'b0,x256 }  )+$signed( { 1'b0,x513 }  )+$signed( { 1'b0,x529 }  )-$signed(11'd108);
assign y384=temp_y[384][11] ==1'b1 ? 5'd0 :  
        temp_y[384][8] ==1'b1 ? 5'd31 : 
        temp_y[384][2]==1'b1 ? temp_y[384][7:3]+1'b1 : temp_y[384][7:3];
assign temp_y[448] = 
+$signed( -{ 2'b0,x0 }<<<3'd1 )+$signed( { 2'b0,x512 } <<<3'd1 )+$signed( -{ 2'b0,x1 }<<<3'd1 )+$signed( { 1'b0,x257 }  )+$signed( { 1'b0,x513 }  )+$signed( -{ 2'b0,x16 }<<<3'd1 )+$signed( { 1'b0,x272 }  )+$signed( { 1'b0,x528 }  )+$signed( -{ 1'b0,x17 } )+$signed(11'd64);
assign y448=temp_y[448][11] ==1'b1 ? 5'd0 :  
        temp_y[448][8] ==1'b1 ? 5'd31 : 
        temp_y[448][2]==1'b1 ? temp_y[448][7:3]+1'b1 : temp_y[448][7:3];
assign temp_y[512] = 
+$signed( -{ 2'b0,x0 }<<<3'd1 )+$signed( -{ 1'b0,x256 } )+$signed( -{ 3'b0,x1 }<<<3'd2)+$signed( { 1'b0,x16 }  )+$signed( { 1'b0,x272 }  )+$signed( { 3'b0,x17 }<<<3'd2 )+$signed(11'd16);
assign y512=temp_y[512][11] ==1'b1 ? 5'd0 :  
        temp_y[512][8] ==1'b1 ? 5'd31 : 
        temp_y[512][2]==1'b1 ? temp_y[512][7:3]+1'b1 : temp_y[512][7:3];
assign temp_y[576] = 
+$signed( { 2'b0,x256 } <<<3'd1 )+$signed( { 2'b0,x512 } <<<3'd1 )+$signed( -{ 1'b0,x1 } )+$signed( -{ 2'b0,x257 }<<<3'd1 )+$signed( -{ 2'b0,x513 }<<<3'd1 )+$signed( { 2'b0,x272 } <<<3'd1 )+$signed( { 1'b0,x528 }  )+$signed( -{ 2'b0,x273 }<<<3'd1 )-$signed(11'd8);
assign y576=temp_y[576][11] ==1'b1 ? 5'd0 :  
        temp_y[576][8] ==1'b1 ? 5'd31 : 
        temp_y[576][2]==1'b1 ? temp_y[576][7:3]+1'b1 : temp_y[576][7:3];
assign temp_y[1] = 
+$signed( -{ 2'b0,x258 }<<<3'd1 )+$signed( -{ 1'b0,x514 } )+$signed( { 1'b0,x3 }  )+$signed( { 1'b0,x259 }  )+$signed( { 1'b0,x515 }  )+$signed( -{ 2'b0,x274 }<<<3'd1 )+$signed( -{ 2'b0,x530 }<<<3'd1 )+$signed( { 2'b0,x275 } <<<3'd1 )+$signed( { 2'b0,x531 } <<<3'd1 )-$signed(11'd16);
assign y1=temp_y[1][11] ==1'b1 ? 5'd0 :  
        temp_y[1][8] ==1'b1 ? 5'd31 : 
        temp_y[1][2]==1'b1 ? temp_y[1][7:3]+1'b1 : temp_y[1][7:3];
assign temp_y[65] = 
+$signed( { 3'b0,x2 }<<<3'd2 )+$signed( -{ 2'b0,x258 }<<<3'd1 )+$signed( -{ 2'b0,x514 }<<<3'd1 )+$signed( { 2'b0,x3 } <<<3'd1 )+$signed( -{ 3'b0,x259 }<<<3'd2)+$signed( { 1'b0,x515 }  )+$signed( -{ 1'b0,x18 } )+$signed( { 1'b0,x530 }  )+$signed( -{ 2'b0,x19 }<<<3'd1 )+$signed( -{ 1'b0,x275 } )+$signed( { 2'b0,x531 } <<<3'd1 )+$signed(11'd24);
assign y65=temp_y[65][11] ==1'b1 ? 5'd0 :  
        temp_y[65][8] ==1'b1 ? 5'd31 : 
        temp_y[65][2]==1'b1 ? temp_y[65][7:3]+1'b1 : temp_y[65][7:3];
assign temp_y[129] = 
+$signed( { 2'b0,x2 } <<<3'd1 )+$signed( { 2'b0,x258 } <<<3'd1 )+$signed( { 1'b0,x514 }  )+$signed( { 2'b0,x3 } <<<3'd1 )+$signed( -{ 1'b0,x259 } )+$signed( { 1'b0,x515 }  )+$signed( -{ 2'b0,x18 }<<<3'd1 )+$signed( -{ 2'b0,x274 }<<<3'd1 )+$signed( -{ 1'b0,x530 } )+$signed( -{ 1'b0,x19 } )+$signed( -{ 1'b0,x275 } )+$signed( -{ 1'b0,x531 } )+$signed(11'd16);
assign y129=temp_y[129][11] ==1'b1 ? 5'd0 :  
        temp_y[129][8] ==1'b1 ? 5'd31 : 
        temp_y[129][2]==1'b1 ? temp_y[129][7:3]+1'b1 : temp_y[129][7:3];
assign temp_y[193] = 
+$signed( { 1'b0,x2 }  )+$signed( -{ 1'b0,x258 } )+$signed( { 1'b0,x3 }  )+$signed( -{ 1'b0,x259 } )+$signed( { 2'b0,x18 } <<<3'd1 )+$signed( -{ 1'b0,x274 } )+$signed( -{ 1'b0,x530 } )+$signed( { 2'b0,x19 } <<<3'd1 )+$signed( -{ 1'b0,x275 } )+$signed( -{ 2'b0,x531 }<<<3'd1 )+$signed(11'd40);
assign y193=temp_y[193][11] ==1'b1 ? 5'd0 :  
        temp_y[193][8] ==1'b1 ? 5'd31 : 
        temp_y[193][2]==1'b1 ? temp_y[193][7:3]+1'b1 : temp_y[193][7:3];
assign temp_y[257] = 
+$signed( -{ 1'b0,x2 } )+$signed( { 2'b0,x258 } <<<3'd1 )+$signed( -{ 1'b0,x514 } )+$signed( -{ 1'b0,x3 } )+$signed( { 2'b0,x259 } <<<3'd1 )+$signed( -{ 2'b0,x515 }<<<3'd1 )+$signed( -{ 1'b0,x18 } )+$signed( { 2'b0,x274 } <<<3'd1 )+$signed( -{ 1'b0,x530 } )+$signed( -{ 2'b0,x19 }<<<3'd1 )+$signed( { 3'b0,x275 }<<<3'd2 )+$signed( -{ 2'b0,x531 }<<<3'd1 )+$signed(11'd32);
assign y257=temp_y[257][11] ==1'b1 ? 5'd0 :  
        temp_y[257][8] ==1'b1 ? 5'd31 : 
        temp_y[257][2]==1'b1 ? temp_y[257][7:3]+1'b1 : temp_y[257][7:3];
assign temp_y[321] = 
+$signed( -{ 1'b0,x2 } )+$signed( -{ 2'b0,x258 }<<<3'd1 )+$signed( -{ 1'b0,x514 } )+$signed( { 1'b0,x3 }  )+$signed( { 2'b0,x259 } <<<3'd1 )+$signed( { 1'b0,x515 }  )+$signed( { 1'b0,x18 }  )+$signed( { 2'b0,x274 } <<<3'd1 )+$signed( { 2'b0,x530 } <<<3'd1 )+$signed( -{ 1'b0,x19 } )+$signed( -{ 2'b0,x275 }<<<3'd1 )+$signed( -{ 1'b0,x531 } )-$signed(11'd68);
assign y321=temp_y[321][11] ==1'b1 ? 5'd0 :  
        temp_y[321][8] ==1'b1 ? 5'd31 : 
        temp_y[321][2]==1'b1 ? temp_y[321][7:3]+1'b1 : temp_y[321][7:3];
assign temp_y[385] = 
+$signed( { 1'b0,x258 }  )+$signed( { 1'b0,x515 }  )+$signed( { 1'b0,x531 }  )-$signed(11'd108);
assign y385=temp_y[385][11] ==1'b1 ? 5'd0 :  
        temp_y[385][8] ==1'b1 ? 5'd31 : 
        temp_y[385][2]==1'b1 ? temp_y[385][7:3]+1'b1 : temp_y[385][7:3];
assign temp_y[449] = 
+$signed( -{ 2'b0,x2 }<<<3'd1 )+$signed( { 2'b0,x514 } <<<3'd1 )+$signed( -{ 2'b0,x3 }<<<3'd1 )+$signed( { 1'b0,x259 }  )+$signed( { 1'b0,x515 }  )+$signed( -{ 2'b0,x18 }<<<3'd1 )+$signed( { 1'b0,x274 }  )+$signed( { 1'b0,x530 }  )+$signed( -{ 1'b0,x19 } )+$signed(11'd64);
assign y449=temp_y[449][11] ==1'b1 ? 5'd0 :  
        temp_y[449][8] ==1'b1 ? 5'd31 : 
        temp_y[449][2]==1'b1 ? temp_y[449][7:3]+1'b1 : temp_y[449][7:3];
assign temp_y[513] = 
+$signed( -{ 2'b0,x2 }<<<3'd1 )+$signed( -{ 1'b0,x258 } )+$signed( -{ 3'b0,x3 }<<<3'd2)+$signed( { 1'b0,x18 }  )+$signed( { 1'b0,x274 }  )+$signed( { 3'b0,x19 }<<<3'd2 )+$signed(11'd16);
assign y513=temp_y[513][11] ==1'b1 ? 5'd0 :  
        temp_y[513][8] ==1'b1 ? 5'd31 : 
        temp_y[513][2]==1'b1 ? temp_y[513][7:3]+1'b1 : temp_y[513][7:3];
assign temp_y[577] = 
+$signed( { 2'b0,x258 } <<<3'd1 )+$signed( { 2'b0,x514 } <<<3'd1 )+$signed( -{ 1'b0,x3 } )+$signed( -{ 2'b0,x259 }<<<3'd1 )+$signed( -{ 2'b0,x515 }<<<3'd1 )+$signed( { 2'b0,x274 } <<<3'd1 )+$signed( { 1'b0,x530 }  )+$signed( -{ 2'b0,x275 }<<<3'd1 )-$signed(11'd8);
assign y577=temp_y[577][11] ==1'b1 ? 5'd0 :  
        temp_y[577][8] ==1'b1 ? 5'd31 : 
        temp_y[577][2]==1'b1 ? temp_y[577][7:3]+1'b1 : temp_y[577][7:3];
assign temp_y[2] = 
+$signed( -{ 2'b0,x260 }<<<3'd1 )+$signed( -{ 1'b0,x516 } )+$signed( { 1'b0,x5 }  )+$signed( { 1'b0,x261 }  )+$signed( { 1'b0,x517 }  )+$signed( -{ 2'b0,x276 }<<<3'd1 )+$signed( -{ 2'b0,x532 }<<<3'd1 )+$signed( { 2'b0,x277 } <<<3'd1 )+$signed( { 2'b0,x533 } <<<3'd1 )-$signed(11'd16);
assign y2=temp_y[2][11] ==1'b1 ? 5'd0 :  
        temp_y[2][8] ==1'b1 ? 5'd31 : 
        temp_y[2][2]==1'b1 ? temp_y[2][7:3]+1'b1 : temp_y[2][7:3];
assign temp_y[66] = 
+$signed( { 3'b0,x4 }<<<3'd2 )+$signed( -{ 2'b0,x260 }<<<3'd1 )+$signed( -{ 2'b0,x516 }<<<3'd1 )+$signed( { 2'b0,x5 } <<<3'd1 )+$signed( -{ 3'b0,x261 }<<<3'd2)+$signed( { 1'b0,x517 }  )+$signed( -{ 1'b0,x20 } )+$signed( { 1'b0,x532 }  )+$signed( -{ 2'b0,x21 }<<<3'd1 )+$signed( -{ 1'b0,x277 } )+$signed( { 2'b0,x533 } <<<3'd1 )+$signed(11'd24);
assign y66=temp_y[66][11] ==1'b1 ? 5'd0 :  
        temp_y[66][8] ==1'b1 ? 5'd31 : 
        temp_y[66][2]==1'b1 ? temp_y[66][7:3]+1'b1 : temp_y[66][7:3];
assign temp_y[130] = 
+$signed( { 2'b0,x4 } <<<3'd1 )+$signed( { 2'b0,x260 } <<<3'd1 )+$signed( { 1'b0,x516 }  )+$signed( { 2'b0,x5 } <<<3'd1 )+$signed( -{ 1'b0,x261 } )+$signed( { 1'b0,x517 }  )+$signed( -{ 2'b0,x20 }<<<3'd1 )+$signed( -{ 2'b0,x276 }<<<3'd1 )+$signed( -{ 1'b0,x532 } )+$signed( -{ 1'b0,x21 } )+$signed( -{ 1'b0,x277 } )+$signed( -{ 1'b0,x533 } )+$signed(11'd16);
assign y130=temp_y[130][11] ==1'b1 ? 5'd0 :  
        temp_y[130][8] ==1'b1 ? 5'd31 : 
        temp_y[130][2]==1'b1 ? temp_y[130][7:3]+1'b1 : temp_y[130][7:3];
assign temp_y[194] = 
+$signed( { 1'b0,x4 }  )+$signed( -{ 1'b0,x260 } )+$signed( { 1'b0,x5 }  )+$signed( -{ 1'b0,x261 } )+$signed( { 2'b0,x20 } <<<3'd1 )+$signed( -{ 1'b0,x276 } )+$signed( -{ 1'b0,x532 } )+$signed( { 2'b0,x21 } <<<3'd1 )+$signed( -{ 1'b0,x277 } )+$signed( -{ 2'b0,x533 }<<<3'd1 )+$signed(11'd40);
assign y194=temp_y[194][11] ==1'b1 ? 5'd0 :  
        temp_y[194][8] ==1'b1 ? 5'd31 : 
        temp_y[194][2]==1'b1 ? temp_y[194][7:3]+1'b1 : temp_y[194][7:3];
assign temp_y[258] = 
+$signed( -{ 1'b0,x4 } )+$signed( { 2'b0,x260 } <<<3'd1 )+$signed( -{ 1'b0,x516 } )+$signed( -{ 1'b0,x5 } )+$signed( { 2'b0,x261 } <<<3'd1 )+$signed( -{ 2'b0,x517 }<<<3'd1 )+$signed( -{ 1'b0,x20 } )+$signed( { 2'b0,x276 } <<<3'd1 )+$signed( -{ 1'b0,x532 } )+$signed( -{ 2'b0,x21 }<<<3'd1 )+$signed( { 3'b0,x277 }<<<3'd2 )+$signed( -{ 2'b0,x533 }<<<3'd1 )+$signed(11'd32);
assign y258=temp_y[258][11] ==1'b1 ? 5'd0 :  
        temp_y[258][8] ==1'b1 ? 5'd31 : 
        temp_y[258][2]==1'b1 ? temp_y[258][7:3]+1'b1 : temp_y[258][7:3];
assign temp_y[322] = 
+$signed( -{ 1'b0,x4 } )+$signed( -{ 2'b0,x260 }<<<3'd1 )+$signed( -{ 1'b0,x516 } )+$signed( { 1'b0,x5 }  )+$signed( { 2'b0,x261 } <<<3'd1 )+$signed( { 1'b0,x517 }  )+$signed( { 1'b0,x20 }  )+$signed( { 2'b0,x276 } <<<3'd1 )+$signed( { 2'b0,x532 } <<<3'd1 )+$signed( -{ 1'b0,x21 } )+$signed( -{ 2'b0,x277 }<<<3'd1 )+$signed( -{ 1'b0,x533 } )-$signed(11'd68);
assign y322=temp_y[322][11] ==1'b1 ? 5'd0 :  
        temp_y[322][8] ==1'b1 ? 5'd31 : 
        temp_y[322][2]==1'b1 ? temp_y[322][7:3]+1'b1 : temp_y[322][7:3];
assign temp_y[386] = 
+$signed( { 1'b0,x260 }  )+$signed( { 1'b0,x517 }  )+$signed( { 1'b0,x533 }  )-$signed(11'd108);
assign y386=temp_y[386][11] ==1'b1 ? 5'd0 :  
        temp_y[386][8] ==1'b1 ? 5'd31 : 
        temp_y[386][2]==1'b1 ? temp_y[386][7:3]+1'b1 : temp_y[386][7:3];
assign temp_y[450] = 
+$signed( -{ 2'b0,x4 }<<<3'd1 )+$signed( { 2'b0,x516 } <<<3'd1 )+$signed( -{ 2'b0,x5 }<<<3'd1 )+$signed( { 1'b0,x261 }  )+$signed( { 1'b0,x517 }  )+$signed( -{ 2'b0,x20 }<<<3'd1 )+$signed( { 1'b0,x276 }  )+$signed( { 1'b0,x532 }  )+$signed( -{ 1'b0,x21 } )+$signed(11'd64);
assign y450=temp_y[450][11] ==1'b1 ? 5'd0 :  
        temp_y[450][8] ==1'b1 ? 5'd31 : 
        temp_y[450][2]==1'b1 ? temp_y[450][7:3]+1'b1 : temp_y[450][7:3];
assign temp_y[514] = 
+$signed( -{ 2'b0,x4 }<<<3'd1 )+$signed( -{ 1'b0,x260 } )+$signed( -{ 3'b0,x5 }<<<3'd2)+$signed( { 1'b0,x20 }  )+$signed( { 1'b0,x276 }  )+$signed( { 3'b0,x21 }<<<3'd2 )+$signed(11'd16);
assign y514=temp_y[514][11] ==1'b1 ? 5'd0 :  
        temp_y[514][8] ==1'b1 ? 5'd31 : 
        temp_y[514][2]==1'b1 ? temp_y[514][7:3]+1'b1 : temp_y[514][7:3];
assign temp_y[578] = 
+$signed( { 2'b0,x260 } <<<3'd1 )+$signed( { 2'b0,x516 } <<<3'd1 )+$signed( -{ 1'b0,x5 } )+$signed( -{ 2'b0,x261 }<<<3'd1 )+$signed( -{ 2'b0,x517 }<<<3'd1 )+$signed( { 2'b0,x276 } <<<3'd1 )+$signed( { 1'b0,x532 }  )+$signed( -{ 2'b0,x277 }<<<3'd1 )-$signed(11'd8);
assign y578=temp_y[578][11] ==1'b1 ? 5'd0 :  
        temp_y[578][8] ==1'b1 ? 5'd31 : 
        temp_y[578][2]==1'b1 ? temp_y[578][7:3]+1'b1 : temp_y[578][7:3];
assign temp_y[3] = 
+$signed( -{ 2'b0,x262 }<<<3'd1 )+$signed( -{ 1'b0,x518 } )+$signed( { 1'b0,x7 }  )+$signed( { 1'b0,x263 }  )+$signed( { 1'b0,x519 }  )+$signed( -{ 2'b0,x278 }<<<3'd1 )+$signed( -{ 2'b0,x534 }<<<3'd1 )+$signed( { 2'b0,x279 } <<<3'd1 )+$signed( { 2'b0,x535 } <<<3'd1 )-$signed(11'd16);
assign y3=temp_y[3][11] ==1'b1 ? 5'd0 :  
        temp_y[3][8] ==1'b1 ? 5'd31 : 
        temp_y[3][2]==1'b1 ? temp_y[3][7:3]+1'b1 : temp_y[3][7:3];
assign temp_y[67] = 
+$signed( { 3'b0,x6 }<<<3'd2 )+$signed( -{ 2'b0,x262 }<<<3'd1 )+$signed( -{ 2'b0,x518 }<<<3'd1 )+$signed( { 2'b0,x7 } <<<3'd1 )+$signed( -{ 3'b0,x263 }<<<3'd2)+$signed( { 1'b0,x519 }  )+$signed( -{ 1'b0,x22 } )+$signed( { 1'b0,x534 }  )+$signed( -{ 2'b0,x23 }<<<3'd1 )+$signed( -{ 1'b0,x279 } )+$signed( { 2'b0,x535 } <<<3'd1 )+$signed(11'd24);
assign y67=temp_y[67][11] ==1'b1 ? 5'd0 :  
        temp_y[67][8] ==1'b1 ? 5'd31 : 
        temp_y[67][2]==1'b1 ? temp_y[67][7:3]+1'b1 : temp_y[67][7:3];
assign temp_y[131] = 
+$signed( { 2'b0,x6 } <<<3'd1 )+$signed( { 2'b0,x262 } <<<3'd1 )+$signed( { 1'b0,x518 }  )+$signed( { 2'b0,x7 } <<<3'd1 )+$signed( -{ 1'b0,x263 } )+$signed( { 1'b0,x519 }  )+$signed( -{ 2'b0,x22 }<<<3'd1 )+$signed( -{ 2'b0,x278 }<<<3'd1 )+$signed( -{ 1'b0,x534 } )+$signed( -{ 1'b0,x23 } )+$signed( -{ 1'b0,x279 } )+$signed( -{ 1'b0,x535 } )+$signed(11'd16);
assign y131=temp_y[131][11] ==1'b1 ? 5'd0 :  
        temp_y[131][8] ==1'b1 ? 5'd31 : 
        temp_y[131][2]==1'b1 ? temp_y[131][7:3]+1'b1 : temp_y[131][7:3];
assign temp_y[195] = 
+$signed( { 1'b0,x6 }  )+$signed( -{ 1'b0,x262 } )+$signed( { 1'b0,x7 }  )+$signed( -{ 1'b0,x263 } )+$signed( { 2'b0,x22 } <<<3'd1 )+$signed( -{ 1'b0,x278 } )+$signed( -{ 1'b0,x534 } )+$signed( { 2'b0,x23 } <<<3'd1 )+$signed( -{ 1'b0,x279 } )+$signed( -{ 2'b0,x535 }<<<3'd1 )+$signed(11'd40);
assign y195=temp_y[195][11] ==1'b1 ? 5'd0 :  
        temp_y[195][8] ==1'b1 ? 5'd31 : 
        temp_y[195][2]==1'b1 ? temp_y[195][7:3]+1'b1 : temp_y[195][7:3];
assign temp_y[259] = 
+$signed( -{ 1'b0,x6 } )+$signed( { 2'b0,x262 } <<<3'd1 )+$signed( -{ 1'b0,x518 } )+$signed( -{ 1'b0,x7 } )+$signed( { 2'b0,x263 } <<<3'd1 )+$signed( -{ 2'b0,x519 }<<<3'd1 )+$signed( -{ 1'b0,x22 } )+$signed( { 2'b0,x278 } <<<3'd1 )+$signed( -{ 1'b0,x534 } )+$signed( -{ 2'b0,x23 }<<<3'd1 )+$signed( { 3'b0,x279 }<<<3'd2 )+$signed( -{ 2'b0,x535 }<<<3'd1 )+$signed(11'd32);
assign y259=temp_y[259][11] ==1'b1 ? 5'd0 :  
        temp_y[259][8] ==1'b1 ? 5'd31 : 
        temp_y[259][2]==1'b1 ? temp_y[259][7:3]+1'b1 : temp_y[259][7:3];
assign temp_y[323] = 
+$signed( -{ 1'b0,x6 } )+$signed( -{ 2'b0,x262 }<<<3'd1 )+$signed( -{ 1'b0,x518 } )+$signed( { 1'b0,x7 }  )+$signed( { 2'b0,x263 } <<<3'd1 )+$signed( { 1'b0,x519 }  )+$signed( { 1'b0,x22 }  )+$signed( { 2'b0,x278 } <<<3'd1 )+$signed( { 2'b0,x534 } <<<3'd1 )+$signed( -{ 1'b0,x23 } )+$signed( -{ 2'b0,x279 }<<<3'd1 )+$signed( -{ 1'b0,x535 } )-$signed(11'd68);
assign y323=temp_y[323][11] ==1'b1 ? 5'd0 :  
        temp_y[323][8] ==1'b1 ? 5'd31 : 
        temp_y[323][2]==1'b1 ? temp_y[323][7:3]+1'b1 : temp_y[323][7:3];
assign temp_y[387] = 
+$signed( { 1'b0,x262 }  )+$signed( { 1'b0,x519 }  )+$signed( { 1'b0,x535 }  )-$signed(11'd108);
assign y387=temp_y[387][11] ==1'b1 ? 5'd0 :  
        temp_y[387][8] ==1'b1 ? 5'd31 : 
        temp_y[387][2]==1'b1 ? temp_y[387][7:3]+1'b1 : temp_y[387][7:3];
assign temp_y[451] = 
+$signed( -{ 2'b0,x6 }<<<3'd1 )+$signed( { 2'b0,x518 } <<<3'd1 )+$signed( -{ 2'b0,x7 }<<<3'd1 )+$signed( { 1'b0,x263 }  )+$signed( { 1'b0,x519 }  )+$signed( -{ 2'b0,x22 }<<<3'd1 )+$signed( { 1'b0,x278 }  )+$signed( { 1'b0,x534 }  )+$signed( -{ 1'b0,x23 } )+$signed(11'd64);
assign y451=temp_y[451][11] ==1'b1 ? 5'd0 :  
        temp_y[451][8] ==1'b1 ? 5'd31 : 
        temp_y[451][2]==1'b1 ? temp_y[451][7:3]+1'b1 : temp_y[451][7:3];
assign temp_y[515] = 
+$signed( -{ 2'b0,x6 }<<<3'd1 )+$signed( -{ 1'b0,x262 } )+$signed( -{ 3'b0,x7 }<<<3'd2)+$signed( { 1'b0,x22 }  )+$signed( { 1'b0,x278 }  )+$signed( { 3'b0,x23 }<<<3'd2 )+$signed(11'd16);
assign y515=temp_y[515][11] ==1'b1 ? 5'd0 :  
        temp_y[515][8] ==1'b1 ? 5'd31 : 
        temp_y[515][2]==1'b1 ? temp_y[515][7:3]+1'b1 : temp_y[515][7:3];
assign temp_y[579] = 
+$signed( { 2'b0,x262 } <<<3'd1 )+$signed( { 2'b0,x518 } <<<3'd1 )+$signed( -{ 1'b0,x7 } )+$signed( -{ 2'b0,x263 }<<<3'd1 )+$signed( -{ 2'b0,x519 }<<<3'd1 )+$signed( { 2'b0,x278 } <<<3'd1 )+$signed( { 1'b0,x534 }  )+$signed( -{ 2'b0,x279 }<<<3'd1 )-$signed(11'd8);
assign y579=temp_y[579][11] ==1'b1 ? 5'd0 :  
        temp_y[579][8] ==1'b1 ? 5'd31 : 
        temp_y[579][2]==1'b1 ? temp_y[579][7:3]+1'b1 : temp_y[579][7:3];
assign temp_y[4] = 
+$signed( -{ 2'b0,x264 }<<<3'd1 )+$signed( -{ 1'b0,x520 } )+$signed( { 1'b0,x9 }  )+$signed( { 1'b0,x265 }  )+$signed( { 1'b0,x521 }  )+$signed( -{ 2'b0,x280 }<<<3'd1 )+$signed( -{ 2'b0,x536 }<<<3'd1 )+$signed( { 2'b0,x281 } <<<3'd1 )+$signed( { 2'b0,x537 } <<<3'd1 )-$signed(11'd16);
assign y4=temp_y[4][11] ==1'b1 ? 5'd0 :  
        temp_y[4][8] ==1'b1 ? 5'd31 : 
        temp_y[4][2]==1'b1 ? temp_y[4][7:3]+1'b1 : temp_y[4][7:3];
assign temp_y[68] = 
+$signed( { 3'b0,x8 }<<<3'd2 )+$signed( -{ 2'b0,x264 }<<<3'd1 )+$signed( -{ 2'b0,x520 }<<<3'd1 )+$signed( { 2'b0,x9 } <<<3'd1 )+$signed( -{ 3'b0,x265 }<<<3'd2)+$signed( { 1'b0,x521 }  )+$signed( -{ 1'b0,x24 } )+$signed( { 1'b0,x536 }  )+$signed( -{ 2'b0,x25 }<<<3'd1 )+$signed( -{ 1'b0,x281 } )+$signed( { 2'b0,x537 } <<<3'd1 )+$signed(11'd24);
assign y68=temp_y[68][11] ==1'b1 ? 5'd0 :  
        temp_y[68][8] ==1'b1 ? 5'd31 : 
        temp_y[68][2]==1'b1 ? temp_y[68][7:3]+1'b1 : temp_y[68][7:3];
assign temp_y[132] = 
+$signed( { 2'b0,x8 } <<<3'd1 )+$signed( { 2'b0,x264 } <<<3'd1 )+$signed( { 1'b0,x520 }  )+$signed( { 2'b0,x9 } <<<3'd1 )+$signed( -{ 1'b0,x265 } )+$signed( { 1'b0,x521 }  )+$signed( -{ 2'b0,x24 }<<<3'd1 )+$signed( -{ 2'b0,x280 }<<<3'd1 )+$signed( -{ 1'b0,x536 } )+$signed( -{ 1'b0,x25 } )+$signed( -{ 1'b0,x281 } )+$signed( -{ 1'b0,x537 } )+$signed(11'd16);
assign y132=temp_y[132][11] ==1'b1 ? 5'd0 :  
        temp_y[132][8] ==1'b1 ? 5'd31 : 
        temp_y[132][2]==1'b1 ? temp_y[132][7:3]+1'b1 : temp_y[132][7:3];
assign temp_y[196] = 
+$signed( { 1'b0,x8 }  )+$signed( -{ 1'b0,x264 } )+$signed( { 1'b0,x9 }  )+$signed( -{ 1'b0,x265 } )+$signed( { 2'b0,x24 } <<<3'd1 )+$signed( -{ 1'b0,x280 } )+$signed( -{ 1'b0,x536 } )+$signed( { 2'b0,x25 } <<<3'd1 )+$signed( -{ 1'b0,x281 } )+$signed( -{ 2'b0,x537 }<<<3'd1 )+$signed(11'd40);
assign y196=temp_y[196][11] ==1'b1 ? 5'd0 :  
        temp_y[196][8] ==1'b1 ? 5'd31 : 
        temp_y[196][2]==1'b1 ? temp_y[196][7:3]+1'b1 : temp_y[196][7:3];
assign temp_y[260] = 
+$signed( -{ 1'b0,x8 } )+$signed( { 2'b0,x264 } <<<3'd1 )+$signed( -{ 1'b0,x520 } )+$signed( -{ 1'b0,x9 } )+$signed( { 2'b0,x265 } <<<3'd1 )+$signed( -{ 2'b0,x521 }<<<3'd1 )+$signed( -{ 1'b0,x24 } )+$signed( { 2'b0,x280 } <<<3'd1 )+$signed( -{ 1'b0,x536 } )+$signed( -{ 2'b0,x25 }<<<3'd1 )+$signed( { 3'b0,x281 }<<<3'd2 )+$signed( -{ 2'b0,x537 }<<<3'd1 )+$signed(11'd32);
assign y260=temp_y[260][11] ==1'b1 ? 5'd0 :  
        temp_y[260][8] ==1'b1 ? 5'd31 : 
        temp_y[260][2]==1'b1 ? temp_y[260][7:3]+1'b1 : temp_y[260][7:3];
assign temp_y[324] = 
+$signed( -{ 1'b0,x8 } )+$signed( -{ 2'b0,x264 }<<<3'd1 )+$signed( -{ 1'b0,x520 } )+$signed( { 1'b0,x9 }  )+$signed( { 2'b0,x265 } <<<3'd1 )+$signed( { 1'b0,x521 }  )+$signed( { 1'b0,x24 }  )+$signed( { 2'b0,x280 } <<<3'd1 )+$signed( { 2'b0,x536 } <<<3'd1 )+$signed( -{ 1'b0,x25 } )+$signed( -{ 2'b0,x281 }<<<3'd1 )+$signed( -{ 1'b0,x537 } )-$signed(11'd68);
assign y324=temp_y[324][11] ==1'b1 ? 5'd0 :  
        temp_y[324][8] ==1'b1 ? 5'd31 : 
        temp_y[324][2]==1'b1 ? temp_y[324][7:3]+1'b1 : temp_y[324][7:3];
assign temp_y[388] = 
+$signed( { 1'b0,x264 }  )+$signed( { 1'b0,x521 }  )+$signed( { 1'b0,x537 }  )-$signed(11'd108);
assign y388=temp_y[388][11] ==1'b1 ? 5'd0 :  
        temp_y[388][8] ==1'b1 ? 5'd31 : 
        temp_y[388][2]==1'b1 ? temp_y[388][7:3]+1'b1 : temp_y[388][7:3];
assign temp_y[452] = 
+$signed( -{ 2'b0,x8 }<<<3'd1 )+$signed( { 2'b0,x520 } <<<3'd1 )+$signed( -{ 2'b0,x9 }<<<3'd1 )+$signed( { 1'b0,x265 }  )+$signed( { 1'b0,x521 }  )+$signed( -{ 2'b0,x24 }<<<3'd1 )+$signed( { 1'b0,x280 }  )+$signed( { 1'b0,x536 }  )+$signed( -{ 1'b0,x25 } )+$signed(11'd64);
assign y452=temp_y[452][11] ==1'b1 ? 5'd0 :  
        temp_y[452][8] ==1'b1 ? 5'd31 : 
        temp_y[452][2]==1'b1 ? temp_y[452][7:3]+1'b1 : temp_y[452][7:3];
assign temp_y[516] = 
+$signed( -{ 2'b0,x8 }<<<3'd1 )+$signed( -{ 1'b0,x264 } )+$signed( -{ 3'b0,x9 }<<<3'd2)+$signed( { 1'b0,x24 }  )+$signed( { 1'b0,x280 }  )+$signed( { 3'b0,x25 }<<<3'd2 )+$signed(11'd16);
assign y516=temp_y[516][11] ==1'b1 ? 5'd0 :  
        temp_y[516][8] ==1'b1 ? 5'd31 : 
        temp_y[516][2]==1'b1 ? temp_y[516][7:3]+1'b1 : temp_y[516][7:3];
assign temp_y[580] = 
+$signed( { 2'b0,x264 } <<<3'd1 )+$signed( { 2'b0,x520 } <<<3'd1 )+$signed( -{ 1'b0,x9 } )+$signed( -{ 2'b0,x265 }<<<3'd1 )+$signed( -{ 2'b0,x521 }<<<3'd1 )+$signed( { 2'b0,x280 } <<<3'd1 )+$signed( { 1'b0,x536 }  )+$signed( -{ 2'b0,x281 }<<<3'd1 )-$signed(11'd8);
assign y580=temp_y[580][11] ==1'b1 ? 5'd0 :  
        temp_y[580][8] ==1'b1 ? 5'd31 : 
        temp_y[580][2]==1'b1 ? temp_y[580][7:3]+1'b1 : temp_y[580][7:3];
assign temp_y[5] = 
+$signed( -{ 2'b0,x266 }<<<3'd1 )+$signed( -{ 1'b0,x522 } )+$signed( { 1'b0,x11 }  )+$signed( { 1'b0,x267 }  )+$signed( { 1'b0,x523 }  )+$signed( -{ 2'b0,x282 }<<<3'd1 )+$signed( -{ 2'b0,x538 }<<<3'd1 )+$signed( { 2'b0,x283 } <<<3'd1 )+$signed( { 2'b0,x539 } <<<3'd1 )-$signed(11'd16);
assign y5=temp_y[5][11] ==1'b1 ? 5'd0 :  
        temp_y[5][8] ==1'b1 ? 5'd31 : 
        temp_y[5][2]==1'b1 ? temp_y[5][7:3]+1'b1 : temp_y[5][7:3];
assign temp_y[69] = 
+$signed( { 3'b0,x10 }<<<3'd2 )+$signed( -{ 2'b0,x266 }<<<3'd1 )+$signed( -{ 2'b0,x522 }<<<3'd1 )+$signed( { 2'b0,x11 } <<<3'd1 )+$signed( -{ 3'b0,x267 }<<<3'd2)+$signed( { 1'b0,x523 }  )+$signed( -{ 1'b0,x26 } )+$signed( { 1'b0,x538 }  )+$signed( -{ 2'b0,x27 }<<<3'd1 )+$signed( -{ 1'b0,x283 } )+$signed( { 2'b0,x539 } <<<3'd1 )+$signed(11'd24);
assign y69=temp_y[69][11] ==1'b1 ? 5'd0 :  
        temp_y[69][8] ==1'b1 ? 5'd31 : 
        temp_y[69][2]==1'b1 ? temp_y[69][7:3]+1'b1 : temp_y[69][7:3];
assign temp_y[133] = 
+$signed( { 2'b0,x10 } <<<3'd1 )+$signed( { 2'b0,x266 } <<<3'd1 )+$signed( { 1'b0,x522 }  )+$signed( { 2'b0,x11 } <<<3'd1 )+$signed( -{ 1'b0,x267 } )+$signed( { 1'b0,x523 }  )+$signed( -{ 2'b0,x26 }<<<3'd1 )+$signed( -{ 2'b0,x282 }<<<3'd1 )+$signed( -{ 1'b0,x538 } )+$signed( -{ 1'b0,x27 } )+$signed( -{ 1'b0,x283 } )+$signed( -{ 1'b0,x539 } )+$signed(11'd16);
assign y133=temp_y[133][11] ==1'b1 ? 5'd0 :  
        temp_y[133][8] ==1'b1 ? 5'd31 : 
        temp_y[133][2]==1'b1 ? temp_y[133][7:3]+1'b1 : temp_y[133][7:3];
assign temp_y[197] = 
+$signed( { 1'b0,x10 }  )+$signed( -{ 1'b0,x266 } )+$signed( { 1'b0,x11 }  )+$signed( -{ 1'b0,x267 } )+$signed( { 2'b0,x26 } <<<3'd1 )+$signed( -{ 1'b0,x282 } )+$signed( -{ 1'b0,x538 } )+$signed( { 2'b0,x27 } <<<3'd1 )+$signed( -{ 1'b0,x283 } )+$signed( -{ 2'b0,x539 }<<<3'd1 )+$signed(11'd40);
assign y197=temp_y[197][11] ==1'b1 ? 5'd0 :  
        temp_y[197][8] ==1'b1 ? 5'd31 : 
        temp_y[197][2]==1'b1 ? temp_y[197][7:3]+1'b1 : temp_y[197][7:3];
assign temp_y[261] = 
+$signed( -{ 1'b0,x10 } )+$signed( { 2'b0,x266 } <<<3'd1 )+$signed( -{ 1'b0,x522 } )+$signed( -{ 1'b0,x11 } )+$signed( { 2'b0,x267 } <<<3'd1 )+$signed( -{ 2'b0,x523 }<<<3'd1 )+$signed( -{ 1'b0,x26 } )+$signed( { 2'b0,x282 } <<<3'd1 )+$signed( -{ 1'b0,x538 } )+$signed( -{ 2'b0,x27 }<<<3'd1 )+$signed( { 3'b0,x283 }<<<3'd2 )+$signed( -{ 2'b0,x539 }<<<3'd1 )+$signed(11'd32);
assign y261=temp_y[261][11] ==1'b1 ? 5'd0 :  
        temp_y[261][8] ==1'b1 ? 5'd31 : 
        temp_y[261][2]==1'b1 ? temp_y[261][7:3]+1'b1 : temp_y[261][7:3];
assign temp_y[325] = 
+$signed( -{ 1'b0,x10 } )+$signed( -{ 2'b0,x266 }<<<3'd1 )+$signed( -{ 1'b0,x522 } )+$signed( { 1'b0,x11 }  )+$signed( { 2'b0,x267 } <<<3'd1 )+$signed( { 1'b0,x523 }  )+$signed( { 1'b0,x26 }  )+$signed( { 2'b0,x282 } <<<3'd1 )+$signed( { 2'b0,x538 } <<<3'd1 )+$signed( -{ 1'b0,x27 } )+$signed( -{ 2'b0,x283 }<<<3'd1 )+$signed( -{ 1'b0,x539 } )-$signed(11'd68);
assign y325=temp_y[325][11] ==1'b1 ? 5'd0 :  
        temp_y[325][8] ==1'b1 ? 5'd31 : 
        temp_y[325][2]==1'b1 ? temp_y[325][7:3]+1'b1 : temp_y[325][7:3];
assign temp_y[389] = 
+$signed( { 1'b0,x266 }  )+$signed( { 1'b0,x523 }  )+$signed( { 1'b0,x539 }  )-$signed(11'd108);
assign y389=temp_y[389][11] ==1'b1 ? 5'd0 :  
        temp_y[389][8] ==1'b1 ? 5'd31 : 
        temp_y[389][2]==1'b1 ? temp_y[389][7:3]+1'b1 : temp_y[389][7:3];
assign temp_y[453] = 
+$signed( -{ 2'b0,x10 }<<<3'd1 )+$signed( { 2'b0,x522 } <<<3'd1 )+$signed( -{ 2'b0,x11 }<<<3'd1 )+$signed( { 1'b0,x267 }  )+$signed( { 1'b0,x523 }  )+$signed( -{ 2'b0,x26 }<<<3'd1 )+$signed( { 1'b0,x282 }  )+$signed( { 1'b0,x538 }  )+$signed( -{ 1'b0,x27 } )+$signed(11'd64);
assign y453=temp_y[453][11] ==1'b1 ? 5'd0 :  
        temp_y[453][8] ==1'b1 ? 5'd31 : 
        temp_y[453][2]==1'b1 ? temp_y[453][7:3]+1'b1 : temp_y[453][7:3];
assign temp_y[517] = 
+$signed( -{ 2'b0,x10 }<<<3'd1 )+$signed( -{ 1'b0,x266 } )+$signed( -{ 3'b0,x11 }<<<3'd2)+$signed( { 1'b0,x26 }  )+$signed( { 1'b0,x282 }  )+$signed( { 3'b0,x27 }<<<3'd2 )+$signed(11'd16);
assign y517=temp_y[517][11] ==1'b1 ? 5'd0 :  
        temp_y[517][8] ==1'b1 ? 5'd31 : 
        temp_y[517][2]==1'b1 ? temp_y[517][7:3]+1'b1 : temp_y[517][7:3];
assign temp_y[581] = 
+$signed( { 2'b0,x266 } <<<3'd1 )+$signed( { 2'b0,x522 } <<<3'd1 )+$signed( -{ 1'b0,x11 } )+$signed( -{ 2'b0,x267 }<<<3'd1 )+$signed( -{ 2'b0,x523 }<<<3'd1 )+$signed( { 2'b0,x282 } <<<3'd1 )+$signed( { 1'b0,x538 }  )+$signed( -{ 2'b0,x283 }<<<3'd1 )-$signed(11'd8);
assign y581=temp_y[581][11] ==1'b1 ? 5'd0 :  
        temp_y[581][8] ==1'b1 ? 5'd31 : 
        temp_y[581][2]==1'b1 ? temp_y[581][7:3]+1'b1 : temp_y[581][7:3];
assign temp_y[6] = 
+$signed( -{ 2'b0,x268 }<<<3'd1 )+$signed( -{ 1'b0,x524 } )+$signed( { 1'b0,x13 }  )+$signed( { 1'b0,x269 }  )+$signed( { 1'b0,x525 }  )+$signed( -{ 2'b0,x284 }<<<3'd1 )+$signed( -{ 2'b0,x540 }<<<3'd1 )+$signed( { 2'b0,x285 } <<<3'd1 )+$signed( { 2'b0,x541 } <<<3'd1 )-$signed(11'd16);
assign y6=temp_y[6][11] ==1'b1 ? 5'd0 :  
        temp_y[6][8] ==1'b1 ? 5'd31 : 
        temp_y[6][2]==1'b1 ? temp_y[6][7:3]+1'b1 : temp_y[6][7:3];
assign temp_y[70] = 
+$signed( { 3'b0,x12 }<<<3'd2 )+$signed( -{ 2'b0,x268 }<<<3'd1 )+$signed( -{ 2'b0,x524 }<<<3'd1 )+$signed( { 2'b0,x13 } <<<3'd1 )+$signed( -{ 3'b0,x269 }<<<3'd2)+$signed( { 1'b0,x525 }  )+$signed( -{ 1'b0,x28 } )+$signed( { 1'b0,x540 }  )+$signed( -{ 2'b0,x29 }<<<3'd1 )+$signed( -{ 1'b0,x285 } )+$signed( { 2'b0,x541 } <<<3'd1 )+$signed(11'd24);
assign y70=temp_y[70][11] ==1'b1 ? 5'd0 :  
        temp_y[70][8] ==1'b1 ? 5'd31 : 
        temp_y[70][2]==1'b1 ? temp_y[70][7:3]+1'b1 : temp_y[70][7:3];
assign temp_y[134] = 
+$signed( { 2'b0,x12 } <<<3'd1 )+$signed( { 2'b0,x268 } <<<3'd1 )+$signed( { 1'b0,x524 }  )+$signed( { 2'b0,x13 } <<<3'd1 )+$signed( -{ 1'b0,x269 } )+$signed( { 1'b0,x525 }  )+$signed( -{ 2'b0,x28 }<<<3'd1 )+$signed( -{ 2'b0,x284 }<<<3'd1 )+$signed( -{ 1'b0,x540 } )+$signed( -{ 1'b0,x29 } )+$signed( -{ 1'b0,x285 } )+$signed( -{ 1'b0,x541 } )+$signed(11'd16);
assign y134=temp_y[134][11] ==1'b1 ? 5'd0 :  
        temp_y[134][8] ==1'b1 ? 5'd31 : 
        temp_y[134][2]==1'b1 ? temp_y[134][7:3]+1'b1 : temp_y[134][7:3];
assign temp_y[198] = 
+$signed( { 1'b0,x12 }  )+$signed( -{ 1'b0,x268 } )+$signed( { 1'b0,x13 }  )+$signed( -{ 1'b0,x269 } )+$signed( { 2'b0,x28 } <<<3'd1 )+$signed( -{ 1'b0,x284 } )+$signed( -{ 1'b0,x540 } )+$signed( { 2'b0,x29 } <<<3'd1 )+$signed( -{ 1'b0,x285 } )+$signed( -{ 2'b0,x541 }<<<3'd1 )+$signed(11'd40);
assign y198=temp_y[198][11] ==1'b1 ? 5'd0 :  
        temp_y[198][8] ==1'b1 ? 5'd31 : 
        temp_y[198][2]==1'b1 ? temp_y[198][7:3]+1'b1 : temp_y[198][7:3];
assign temp_y[262] = 
+$signed( -{ 1'b0,x12 } )+$signed( { 2'b0,x268 } <<<3'd1 )+$signed( -{ 1'b0,x524 } )+$signed( -{ 1'b0,x13 } )+$signed( { 2'b0,x269 } <<<3'd1 )+$signed( -{ 2'b0,x525 }<<<3'd1 )+$signed( -{ 1'b0,x28 } )+$signed( { 2'b0,x284 } <<<3'd1 )+$signed( -{ 1'b0,x540 } )+$signed( -{ 2'b0,x29 }<<<3'd1 )+$signed( { 3'b0,x285 }<<<3'd2 )+$signed( -{ 2'b0,x541 }<<<3'd1 )+$signed(11'd32);
assign y262=temp_y[262][11] ==1'b1 ? 5'd0 :  
        temp_y[262][8] ==1'b1 ? 5'd31 : 
        temp_y[262][2]==1'b1 ? temp_y[262][7:3]+1'b1 : temp_y[262][7:3];
assign temp_y[326] = 
+$signed( -{ 1'b0,x12 } )+$signed( -{ 2'b0,x268 }<<<3'd1 )+$signed( -{ 1'b0,x524 } )+$signed( { 1'b0,x13 }  )+$signed( { 2'b0,x269 } <<<3'd1 )+$signed( { 1'b0,x525 }  )+$signed( { 1'b0,x28 }  )+$signed( { 2'b0,x284 } <<<3'd1 )+$signed( { 2'b0,x540 } <<<3'd1 )+$signed( -{ 1'b0,x29 } )+$signed( -{ 2'b0,x285 }<<<3'd1 )+$signed( -{ 1'b0,x541 } )-$signed(11'd68);
assign y326=temp_y[326][11] ==1'b1 ? 5'd0 :  
        temp_y[326][8] ==1'b1 ? 5'd31 : 
        temp_y[326][2]==1'b1 ? temp_y[326][7:3]+1'b1 : temp_y[326][7:3];
assign temp_y[390] = 
+$signed( { 1'b0,x268 }  )+$signed( { 1'b0,x525 }  )+$signed( { 1'b0,x541 }  )-$signed(11'd108);
assign y390=temp_y[390][11] ==1'b1 ? 5'd0 :  
        temp_y[390][8] ==1'b1 ? 5'd31 : 
        temp_y[390][2]==1'b1 ? temp_y[390][7:3]+1'b1 : temp_y[390][7:3];
assign temp_y[454] = 
+$signed( -{ 2'b0,x12 }<<<3'd1 )+$signed( { 2'b0,x524 } <<<3'd1 )+$signed( -{ 2'b0,x13 }<<<3'd1 )+$signed( { 1'b0,x269 }  )+$signed( { 1'b0,x525 }  )+$signed( -{ 2'b0,x28 }<<<3'd1 )+$signed( { 1'b0,x284 }  )+$signed( { 1'b0,x540 }  )+$signed( -{ 1'b0,x29 } )+$signed(11'd64);
assign y454=temp_y[454][11] ==1'b1 ? 5'd0 :  
        temp_y[454][8] ==1'b1 ? 5'd31 : 
        temp_y[454][2]==1'b1 ? temp_y[454][7:3]+1'b1 : temp_y[454][7:3];
assign temp_y[518] = 
+$signed( -{ 2'b0,x12 }<<<3'd1 )+$signed( -{ 1'b0,x268 } )+$signed( -{ 3'b0,x13 }<<<3'd2)+$signed( { 1'b0,x28 }  )+$signed( { 1'b0,x284 }  )+$signed( { 3'b0,x29 }<<<3'd2 )+$signed(11'd16);
assign y518=temp_y[518][11] ==1'b1 ? 5'd0 :  
        temp_y[518][8] ==1'b1 ? 5'd31 : 
        temp_y[518][2]==1'b1 ? temp_y[518][7:3]+1'b1 : temp_y[518][7:3];
assign temp_y[582] = 
+$signed( { 2'b0,x268 } <<<3'd1 )+$signed( { 2'b0,x524 } <<<3'd1 )+$signed( -{ 1'b0,x13 } )+$signed( -{ 2'b0,x269 }<<<3'd1 )+$signed( -{ 2'b0,x525 }<<<3'd1 )+$signed( { 2'b0,x284 } <<<3'd1 )+$signed( { 1'b0,x540 }  )+$signed( -{ 2'b0,x285 }<<<3'd1 )-$signed(11'd8);
assign y582=temp_y[582][11] ==1'b1 ? 5'd0 :  
        temp_y[582][8] ==1'b1 ? 5'd31 : 
        temp_y[582][2]==1'b1 ? temp_y[582][7:3]+1'b1 : temp_y[582][7:3];
assign temp_y[7] = 
+$signed( -{ 2'b0,x270 }<<<3'd1 )+$signed( -{ 1'b0,x526 } )+$signed( { 1'b0,x15 }  )+$signed( { 1'b0,x271 }  )+$signed( { 1'b0,x527 }  )+$signed( -{ 2'b0,x286 }<<<3'd1 )+$signed( -{ 2'b0,x542 }<<<3'd1 )+$signed( { 2'b0,x287 } <<<3'd1 )+$signed( { 2'b0,x543 } <<<3'd1 )-$signed(11'd16);
assign y7=temp_y[7][11] ==1'b1 ? 5'd0 :  
        temp_y[7][8] ==1'b1 ? 5'd31 : 
        temp_y[7][2]==1'b1 ? temp_y[7][7:3]+1'b1 : temp_y[7][7:3];
assign temp_y[71] = 
+$signed( { 3'b0,x14 }<<<3'd2 )+$signed( -{ 2'b0,x270 }<<<3'd1 )+$signed( -{ 2'b0,x526 }<<<3'd1 )+$signed( { 2'b0,x15 } <<<3'd1 )+$signed( -{ 3'b0,x271 }<<<3'd2)+$signed( { 1'b0,x527 }  )+$signed( -{ 1'b0,x30 } )+$signed( { 1'b0,x542 }  )+$signed( -{ 2'b0,x31 }<<<3'd1 )+$signed( -{ 1'b0,x287 } )+$signed( { 2'b0,x543 } <<<3'd1 )+$signed(11'd24);
assign y71=temp_y[71][11] ==1'b1 ? 5'd0 :  
        temp_y[71][8] ==1'b1 ? 5'd31 : 
        temp_y[71][2]==1'b1 ? temp_y[71][7:3]+1'b1 : temp_y[71][7:3];
assign temp_y[135] = 
+$signed( { 2'b0,x14 } <<<3'd1 )+$signed( { 2'b0,x270 } <<<3'd1 )+$signed( { 1'b0,x526 }  )+$signed( { 2'b0,x15 } <<<3'd1 )+$signed( -{ 1'b0,x271 } )+$signed( { 1'b0,x527 }  )+$signed( -{ 2'b0,x30 }<<<3'd1 )+$signed( -{ 2'b0,x286 }<<<3'd1 )+$signed( -{ 1'b0,x542 } )+$signed( -{ 1'b0,x31 } )+$signed( -{ 1'b0,x287 } )+$signed( -{ 1'b0,x543 } )+$signed(11'd16);
assign y135=temp_y[135][11] ==1'b1 ? 5'd0 :  
        temp_y[135][8] ==1'b1 ? 5'd31 : 
        temp_y[135][2]==1'b1 ? temp_y[135][7:3]+1'b1 : temp_y[135][7:3];
assign temp_y[199] = 
+$signed( { 1'b0,x14 }  )+$signed( -{ 1'b0,x270 } )+$signed( { 1'b0,x15 }  )+$signed( -{ 1'b0,x271 } )+$signed( { 2'b0,x30 } <<<3'd1 )+$signed( -{ 1'b0,x286 } )+$signed( -{ 1'b0,x542 } )+$signed( { 2'b0,x31 } <<<3'd1 )+$signed( -{ 1'b0,x287 } )+$signed( -{ 2'b0,x543 }<<<3'd1 )+$signed(11'd40);
assign y199=temp_y[199][11] ==1'b1 ? 5'd0 :  
        temp_y[199][8] ==1'b1 ? 5'd31 : 
        temp_y[199][2]==1'b1 ? temp_y[199][7:3]+1'b1 : temp_y[199][7:3];
assign temp_y[263] = 
+$signed( -{ 1'b0,x14 } )+$signed( { 2'b0,x270 } <<<3'd1 )+$signed( -{ 1'b0,x526 } )+$signed( -{ 1'b0,x15 } )+$signed( { 2'b0,x271 } <<<3'd1 )+$signed( -{ 2'b0,x527 }<<<3'd1 )+$signed( -{ 1'b0,x30 } )+$signed( { 2'b0,x286 } <<<3'd1 )+$signed( -{ 1'b0,x542 } )+$signed( -{ 2'b0,x31 }<<<3'd1 )+$signed( { 3'b0,x287 }<<<3'd2 )+$signed( -{ 2'b0,x543 }<<<3'd1 )+$signed(11'd32);
assign y263=temp_y[263][11] ==1'b1 ? 5'd0 :  
        temp_y[263][8] ==1'b1 ? 5'd31 : 
        temp_y[263][2]==1'b1 ? temp_y[263][7:3]+1'b1 : temp_y[263][7:3];
assign temp_y[327] = 
+$signed( -{ 1'b0,x14 } )+$signed( -{ 2'b0,x270 }<<<3'd1 )+$signed( -{ 1'b0,x526 } )+$signed( { 1'b0,x15 }  )+$signed( { 2'b0,x271 } <<<3'd1 )+$signed( { 1'b0,x527 }  )+$signed( { 1'b0,x30 }  )+$signed( { 2'b0,x286 } <<<3'd1 )+$signed( { 2'b0,x542 } <<<3'd1 )+$signed( -{ 1'b0,x31 } )+$signed( -{ 2'b0,x287 }<<<3'd1 )+$signed( -{ 1'b0,x543 } )-$signed(11'd68);
assign y327=temp_y[327][11] ==1'b1 ? 5'd0 :  
        temp_y[327][8] ==1'b1 ? 5'd31 : 
        temp_y[327][2]==1'b1 ? temp_y[327][7:3]+1'b1 : temp_y[327][7:3];
assign temp_y[391] = 
+$signed( { 1'b0,x270 }  )+$signed( { 1'b0,x527 }  )+$signed( { 1'b0,x543 }  )-$signed(11'd108);
assign y391=temp_y[391][11] ==1'b1 ? 5'd0 :  
        temp_y[391][8] ==1'b1 ? 5'd31 : 
        temp_y[391][2]==1'b1 ? temp_y[391][7:3]+1'b1 : temp_y[391][7:3];
assign temp_y[455] = 
+$signed( -{ 2'b0,x14 }<<<3'd1 )+$signed( { 2'b0,x526 } <<<3'd1 )+$signed( -{ 2'b0,x15 }<<<3'd1 )+$signed( { 1'b0,x271 }  )+$signed( { 1'b0,x527 }  )+$signed( -{ 2'b0,x30 }<<<3'd1 )+$signed( { 1'b0,x286 }  )+$signed( { 1'b0,x542 }  )+$signed( -{ 1'b0,x31 } )+$signed(11'd64);
assign y455=temp_y[455][11] ==1'b1 ? 5'd0 :  
        temp_y[455][8] ==1'b1 ? 5'd31 : 
        temp_y[455][2]==1'b1 ? temp_y[455][7:3]+1'b1 : temp_y[455][7:3];
assign temp_y[519] = 
+$signed( -{ 2'b0,x14 }<<<3'd1 )+$signed( -{ 1'b0,x270 } )+$signed( -{ 3'b0,x15 }<<<3'd2)+$signed( { 1'b0,x30 }  )+$signed( { 1'b0,x286 }  )+$signed( { 3'b0,x31 }<<<3'd2 )+$signed(11'd16);
assign y519=temp_y[519][11] ==1'b1 ? 5'd0 :  
        temp_y[519][8] ==1'b1 ? 5'd31 : 
        temp_y[519][2]==1'b1 ? temp_y[519][7:3]+1'b1 : temp_y[519][7:3];
assign temp_y[583] = 
+$signed( { 2'b0,x270 } <<<3'd1 )+$signed( { 2'b0,x526 } <<<3'd1 )+$signed( -{ 1'b0,x15 } )+$signed( -{ 2'b0,x271 }<<<3'd1 )+$signed( -{ 2'b0,x527 }<<<3'd1 )+$signed( { 2'b0,x286 } <<<3'd1 )+$signed( { 1'b0,x542 }  )+$signed( -{ 2'b0,x287 }<<<3'd1 )-$signed(11'd8);
assign y583=temp_y[583][11] ==1'b1 ? 5'd0 :  
        temp_y[583][8] ==1'b1 ? 5'd31 : 
        temp_y[583][2]==1'b1 ? temp_y[583][7:3]+1'b1 : temp_y[583][7:3];
assign temp_y[8] = 
+$signed( -{ 2'b0,x288 }<<<3'd1 )+$signed( -{ 1'b0,x544 } )+$signed( { 1'b0,x33 }  )+$signed( { 1'b0,x289 }  )+$signed( { 1'b0,x545 }  )+$signed( -{ 2'b0,x304 }<<<3'd1 )+$signed( -{ 2'b0,x560 }<<<3'd1 )+$signed( { 2'b0,x305 } <<<3'd1 )+$signed( { 2'b0,x561 } <<<3'd1 )-$signed(11'd16);
assign y8=temp_y[8][11] ==1'b1 ? 5'd0 :  
        temp_y[8][8] ==1'b1 ? 5'd31 : 
        temp_y[8][2]==1'b1 ? temp_y[8][7:3]+1'b1 : temp_y[8][7:3];
assign temp_y[72] = 
+$signed( { 3'b0,x32 }<<<3'd2 )+$signed( -{ 2'b0,x288 }<<<3'd1 )+$signed( -{ 2'b0,x544 }<<<3'd1 )+$signed( { 2'b0,x33 } <<<3'd1 )+$signed( -{ 3'b0,x289 }<<<3'd2)+$signed( { 1'b0,x545 }  )+$signed( -{ 1'b0,x48 } )+$signed( { 1'b0,x560 }  )+$signed( -{ 2'b0,x49 }<<<3'd1 )+$signed( -{ 1'b0,x305 } )+$signed( { 2'b0,x561 } <<<3'd1 )+$signed(11'd24);
assign y72=temp_y[72][11] ==1'b1 ? 5'd0 :  
        temp_y[72][8] ==1'b1 ? 5'd31 : 
        temp_y[72][2]==1'b1 ? temp_y[72][7:3]+1'b1 : temp_y[72][7:3];
assign temp_y[136] = 
+$signed( { 2'b0,x32 } <<<3'd1 )+$signed( { 2'b0,x288 } <<<3'd1 )+$signed( { 1'b0,x544 }  )+$signed( { 2'b0,x33 } <<<3'd1 )+$signed( -{ 1'b0,x289 } )+$signed( { 1'b0,x545 }  )+$signed( -{ 2'b0,x48 }<<<3'd1 )+$signed( -{ 2'b0,x304 }<<<3'd1 )+$signed( -{ 1'b0,x560 } )+$signed( -{ 1'b0,x49 } )+$signed( -{ 1'b0,x305 } )+$signed( -{ 1'b0,x561 } )+$signed(11'd16);
assign y136=temp_y[136][11] ==1'b1 ? 5'd0 :  
        temp_y[136][8] ==1'b1 ? 5'd31 : 
        temp_y[136][2]==1'b1 ? temp_y[136][7:3]+1'b1 : temp_y[136][7:3];
assign temp_y[200] = 
+$signed( { 1'b0,x32 }  )+$signed( -{ 1'b0,x288 } )+$signed( { 1'b0,x33 }  )+$signed( -{ 1'b0,x289 } )+$signed( { 2'b0,x48 } <<<3'd1 )+$signed( -{ 1'b0,x304 } )+$signed( -{ 1'b0,x560 } )+$signed( { 2'b0,x49 } <<<3'd1 )+$signed( -{ 1'b0,x305 } )+$signed( -{ 2'b0,x561 }<<<3'd1 )+$signed(11'd40);
assign y200=temp_y[200][11] ==1'b1 ? 5'd0 :  
        temp_y[200][8] ==1'b1 ? 5'd31 : 
        temp_y[200][2]==1'b1 ? temp_y[200][7:3]+1'b1 : temp_y[200][7:3];
assign temp_y[264] = 
+$signed( -{ 1'b0,x32 } )+$signed( { 2'b0,x288 } <<<3'd1 )+$signed( -{ 1'b0,x544 } )+$signed( -{ 1'b0,x33 } )+$signed( { 2'b0,x289 } <<<3'd1 )+$signed( -{ 2'b0,x545 }<<<3'd1 )+$signed( -{ 1'b0,x48 } )+$signed( { 2'b0,x304 } <<<3'd1 )+$signed( -{ 1'b0,x560 } )+$signed( -{ 2'b0,x49 }<<<3'd1 )+$signed( { 3'b0,x305 }<<<3'd2 )+$signed( -{ 2'b0,x561 }<<<3'd1 )+$signed(11'd32);
assign y264=temp_y[264][11] ==1'b1 ? 5'd0 :  
        temp_y[264][8] ==1'b1 ? 5'd31 : 
        temp_y[264][2]==1'b1 ? temp_y[264][7:3]+1'b1 : temp_y[264][7:3];
assign temp_y[328] = 
+$signed( -{ 1'b0,x32 } )+$signed( -{ 2'b0,x288 }<<<3'd1 )+$signed( -{ 1'b0,x544 } )+$signed( { 1'b0,x33 }  )+$signed( { 2'b0,x289 } <<<3'd1 )+$signed( { 1'b0,x545 }  )+$signed( { 1'b0,x48 }  )+$signed( { 2'b0,x304 } <<<3'd1 )+$signed( { 2'b0,x560 } <<<3'd1 )+$signed( -{ 1'b0,x49 } )+$signed( -{ 2'b0,x305 }<<<3'd1 )+$signed( -{ 1'b0,x561 } )-$signed(11'd68);
assign y328=temp_y[328][11] ==1'b1 ? 5'd0 :  
        temp_y[328][8] ==1'b1 ? 5'd31 : 
        temp_y[328][2]==1'b1 ? temp_y[328][7:3]+1'b1 : temp_y[328][7:3];
assign temp_y[392] = 
+$signed( { 1'b0,x288 }  )+$signed( { 1'b0,x545 }  )+$signed( { 1'b0,x561 }  )-$signed(11'd108);
assign y392=temp_y[392][11] ==1'b1 ? 5'd0 :  
        temp_y[392][8] ==1'b1 ? 5'd31 : 
        temp_y[392][2]==1'b1 ? temp_y[392][7:3]+1'b1 : temp_y[392][7:3];
assign temp_y[456] = 
+$signed( -{ 2'b0,x32 }<<<3'd1 )+$signed( { 2'b0,x544 } <<<3'd1 )+$signed( -{ 2'b0,x33 }<<<3'd1 )+$signed( { 1'b0,x289 }  )+$signed( { 1'b0,x545 }  )+$signed( -{ 2'b0,x48 }<<<3'd1 )+$signed( { 1'b0,x304 }  )+$signed( { 1'b0,x560 }  )+$signed( -{ 1'b0,x49 } )+$signed(11'd64);
assign y456=temp_y[456][11] ==1'b1 ? 5'd0 :  
        temp_y[456][8] ==1'b1 ? 5'd31 : 
        temp_y[456][2]==1'b1 ? temp_y[456][7:3]+1'b1 : temp_y[456][7:3];
assign temp_y[520] = 
+$signed( -{ 2'b0,x32 }<<<3'd1 )+$signed( -{ 1'b0,x288 } )+$signed( -{ 3'b0,x33 }<<<3'd2)+$signed( { 1'b0,x48 }  )+$signed( { 1'b0,x304 }  )+$signed( { 3'b0,x49 }<<<3'd2 )+$signed(11'd16);
assign y520=temp_y[520][11] ==1'b1 ? 5'd0 :  
        temp_y[520][8] ==1'b1 ? 5'd31 : 
        temp_y[520][2]==1'b1 ? temp_y[520][7:3]+1'b1 : temp_y[520][7:3];
assign temp_y[584] = 
+$signed( { 2'b0,x288 } <<<3'd1 )+$signed( { 2'b0,x544 } <<<3'd1 )+$signed( -{ 1'b0,x33 } )+$signed( -{ 2'b0,x289 }<<<3'd1 )+$signed( -{ 2'b0,x545 }<<<3'd1 )+$signed( { 2'b0,x304 } <<<3'd1 )+$signed( { 1'b0,x560 }  )+$signed( -{ 2'b0,x305 }<<<3'd1 )-$signed(11'd8);
assign y584=temp_y[584][11] ==1'b1 ? 5'd0 :  
        temp_y[584][8] ==1'b1 ? 5'd31 : 
        temp_y[584][2]==1'b1 ? temp_y[584][7:3]+1'b1 : temp_y[584][7:3];
assign temp_y[9] = 
+$signed( -{ 2'b0,x290 }<<<3'd1 )+$signed( -{ 1'b0,x546 } )+$signed( { 1'b0,x35 }  )+$signed( { 1'b0,x291 }  )+$signed( { 1'b0,x547 }  )+$signed( -{ 2'b0,x306 }<<<3'd1 )+$signed( -{ 2'b0,x562 }<<<3'd1 )+$signed( { 2'b0,x307 } <<<3'd1 )+$signed( { 2'b0,x563 } <<<3'd1 )-$signed(11'd16);
assign y9=temp_y[9][11] ==1'b1 ? 5'd0 :  
        temp_y[9][8] ==1'b1 ? 5'd31 : 
        temp_y[9][2]==1'b1 ? temp_y[9][7:3]+1'b1 : temp_y[9][7:3];
assign temp_y[73] = 
+$signed( { 3'b0,x34 }<<<3'd2 )+$signed( -{ 2'b0,x290 }<<<3'd1 )+$signed( -{ 2'b0,x546 }<<<3'd1 )+$signed( { 2'b0,x35 } <<<3'd1 )+$signed( -{ 3'b0,x291 }<<<3'd2)+$signed( { 1'b0,x547 }  )+$signed( -{ 1'b0,x50 } )+$signed( { 1'b0,x562 }  )+$signed( -{ 2'b0,x51 }<<<3'd1 )+$signed( -{ 1'b0,x307 } )+$signed( { 2'b0,x563 } <<<3'd1 )+$signed(11'd24);
assign y73=temp_y[73][11] ==1'b1 ? 5'd0 :  
        temp_y[73][8] ==1'b1 ? 5'd31 : 
        temp_y[73][2]==1'b1 ? temp_y[73][7:3]+1'b1 : temp_y[73][7:3];
assign temp_y[137] = 
+$signed( { 2'b0,x34 } <<<3'd1 )+$signed( { 2'b0,x290 } <<<3'd1 )+$signed( { 1'b0,x546 }  )+$signed( { 2'b0,x35 } <<<3'd1 )+$signed( -{ 1'b0,x291 } )+$signed( { 1'b0,x547 }  )+$signed( -{ 2'b0,x50 }<<<3'd1 )+$signed( -{ 2'b0,x306 }<<<3'd1 )+$signed( -{ 1'b0,x562 } )+$signed( -{ 1'b0,x51 } )+$signed( -{ 1'b0,x307 } )+$signed( -{ 1'b0,x563 } )+$signed(11'd16);
assign y137=temp_y[137][11] ==1'b1 ? 5'd0 :  
        temp_y[137][8] ==1'b1 ? 5'd31 : 
        temp_y[137][2]==1'b1 ? temp_y[137][7:3]+1'b1 : temp_y[137][7:3];
assign temp_y[201] = 
+$signed( { 1'b0,x34 }  )+$signed( -{ 1'b0,x290 } )+$signed( { 1'b0,x35 }  )+$signed( -{ 1'b0,x291 } )+$signed( { 2'b0,x50 } <<<3'd1 )+$signed( -{ 1'b0,x306 } )+$signed( -{ 1'b0,x562 } )+$signed( { 2'b0,x51 } <<<3'd1 )+$signed( -{ 1'b0,x307 } )+$signed( -{ 2'b0,x563 }<<<3'd1 )+$signed(11'd40);
assign y201=temp_y[201][11] ==1'b1 ? 5'd0 :  
        temp_y[201][8] ==1'b1 ? 5'd31 : 
        temp_y[201][2]==1'b1 ? temp_y[201][7:3]+1'b1 : temp_y[201][7:3];
assign temp_y[265] = 
+$signed( -{ 1'b0,x34 } )+$signed( { 2'b0,x290 } <<<3'd1 )+$signed( -{ 1'b0,x546 } )+$signed( -{ 1'b0,x35 } )+$signed( { 2'b0,x291 } <<<3'd1 )+$signed( -{ 2'b0,x547 }<<<3'd1 )+$signed( -{ 1'b0,x50 } )+$signed( { 2'b0,x306 } <<<3'd1 )+$signed( -{ 1'b0,x562 } )+$signed( -{ 2'b0,x51 }<<<3'd1 )+$signed( { 3'b0,x307 }<<<3'd2 )+$signed( -{ 2'b0,x563 }<<<3'd1 )+$signed(11'd32);
assign y265=temp_y[265][11] ==1'b1 ? 5'd0 :  
        temp_y[265][8] ==1'b1 ? 5'd31 : 
        temp_y[265][2]==1'b1 ? temp_y[265][7:3]+1'b1 : temp_y[265][7:3];
assign temp_y[329] = 
+$signed( -{ 1'b0,x34 } )+$signed( -{ 2'b0,x290 }<<<3'd1 )+$signed( -{ 1'b0,x546 } )+$signed( { 1'b0,x35 }  )+$signed( { 2'b0,x291 } <<<3'd1 )+$signed( { 1'b0,x547 }  )+$signed( { 1'b0,x50 }  )+$signed( { 2'b0,x306 } <<<3'd1 )+$signed( { 2'b0,x562 } <<<3'd1 )+$signed( -{ 1'b0,x51 } )+$signed( -{ 2'b0,x307 }<<<3'd1 )+$signed( -{ 1'b0,x563 } )-$signed(11'd68);
assign y329=temp_y[329][11] ==1'b1 ? 5'd0 :  
        temp_y[329][8] ==1'b1 ? 5'd31 : 
        temp_y[329][2]==1'b1 ? temp_y[329][7:3]+1'b1 : temp_y[329][7:3];
assign temp_y[393] = 
+$signed( { 1'b0,x290 }  )+$signed( { 1'b0,x547 }  )+$signed( { 1'b0,x563 }  )-$signed(11'd108);
assign y393=temp_y[393][11] ==1'b1 ? 5'd0 :  
        temp_y[393][8] ==1'b1 ? 5'd31 : 
        temp_y[393][2]==1'b1 ? temp_y[393][7:3]+1'b1 : temp_y[393][7:3];
assign temp_y[457] = 
+$signed( -{ 2'b0,x34 }<<<3'd1 )+$signed( { 2'b0,x546 } <<<3'd1 )+$signed( -{ 2'b0,x35 }<<<3'd1 )+$signed( { 1'b0,x291 }  )+$signed( { 1'b0,x547 }  )+$signed( -{ 2'b0,x50 }<<<3'd1 )+$signed( { 1'b0,x306 }  )+$signed( { 1'b0,x562 }  )+$signed( -{ 1'b0,x51 } )+$signed(11'd64);
assign y457=temp_y[457][11] ==1'b1 ? 5'd0 :  
        temp_y[457][8] ==1'b1 ? 5'd31 : 
        temp_y[457][2]==1'b1 ? temp_y[457][7:3]+1'b1 : temp_y[457][7:3];
assign temp_y[521] = 
+$signed( -{ 2'b0,x34 }<<<3'd1 )+$signed( -{ 1'b0,x290 } )+$signed( -{ 3'b0,x35 }<<<3'd2)+$signed( { 1'b0,x50 }  )+$signed( { 1'b0,x306 }  )+$signed( { 3'b0,x51 }<<<3'd2 )+$signed(11'd16);
assign y521=temp_y[521][11] ==1'b1 ? 5'd0 :  
        temp_y[521][8] ==1'b1 ? 5'd31 : 
        temp_y[521][2]==1'b1 ? temp_y[521][7:3]+1'b1 : temp_y[521][7:3];
assign temp_y[585] = 
+$signed( { 2'b0,x290 } <<<3'd1 )+$signed( { 2'b0,x546 } <<<3'd1 )+$signed( -{ 1'b0,x35 } )+$signed( -{ 2'b0,x291 }<<<3'd1 )+$signed( -{ 2'b0,x547 }<<<3'd1 )+$signed( { 2'b0,x306 } <<<3'd1 )+$signed( { 1'b0,x562 }  )+$signed( -{ 2'b0,x307 }<<<3'd1 )-$signed(11'd8);
assign y585=temp_y[585][11] ==1'b1 ? 5'd0 :  
        temp_y[585][8] ==1'b1 ? 5'd31 : 
        temp_y[585][2]==1'b1 ? temp_y[585][7:3]+1'b1 : temp_y[585][7:3];
assign temp_y[10] = 
+$signed( -{ 2'b0,x292 }<<<3'd1 )+$signed( -{ 1'b0,x548 } )+$signed( { 1'b0,x37 }  )+$signed( { 1'b0,x293 }  )+$signed( { 1'b0,x549 }  )+$signed( -{ 2'b0,x308 }<<<3'd1 )+$signed( -{ 2'b0,x564 }<<<3'd1 )+$signed( { 2'b0,x309 } <<<3'd1 )+$signed( { 2'b0,x565 } <<<3'd1 )-$signed(11'd16);
assign y10=temp_y[10][11] ==1'b1 ? 5'd0 :  
        temp_y[10][8] ==1'b1 ? 5'd31 : 
        temp_y[10][2]==1'b1 ? temp_y[10][7:3]+1'b1 : temp_y[10][7:3];
assign temp_y[74] = 
+$signed( { 3'b0,x36 }<<<3'd2 )+$signed( -{ 2'b0,x292 }<<<3'd1 )+$signed( -{ 2'b0,x548 }<<<3'd1 )+$signed( { 2'b0,x37 } <<<3'd1 )+$signed( -{ 3'b0,x293 }<<<3'd2)+$signed( { 1'b0,x549 }  )+$signed( -{ 1'b0,x52 } )+$signed( { 1'b0,x564 }  )+$signed( -{ 2'b0,x53 }<<<3'd1 )+$signed( -{ 1'b0,x309 } )+$signed( { 2'b0,x565 } <<<3'd1 )+$signed(11'd24);
assign y74=temp_y[74][11] ==1'b1 ? 5'd0 :  
        temp_y[74][8] ==1'b1 ? 5'd31 : 
        temp_y[74][2]==1'b1 ? temp_y[74][7:3]+1'b1 : temp_y[74][7:3];
assign temp_y[138] = 
+$signed( { 2'b0,x36 } <<<3'd1 )+$signed( { 2'b0,x292 } <<<3'd1 )+$signed( { 1'b0,x548 }  )+$signed( { 2'b0,x37 } <<<3'd1 )+$signed( -{ 1'b0,x293 } )+$signed( { 1'b0,x549 }  )+$signed( -{ 2'b0,x52 }<<<3'd1 )+$signed( -{ 2'b0,x308 }<<<3'd1 )+$signed( -{ 1'b0,x564 } )+$signed( -{ 1'b0,x53 } )+$signed( -{ 1'b0,x309 } )+$signed( -{ 1'b0,x565 } )+$signed(11'd16);
assign y138=temp_y[138][11] ==1'b1 ? 5'd0 :  
        temp_y[138][8] ==1'b1 ? 5'd31 : 
        temp_y[138][2]==1'b1 ? temp_y[138][7:3]+1'b1 : temp_y[138][7:3];
assign temp_y[202] = 
+$signed( { 1'b0,x36 }  )+$signed( -{ 1'b0,x292 } )+$signed( { 1'b0,x37 }  )+$signed( -{ 1'b0,x293 } )+$signed( { 2'b0,x52 } <<<3'd1 )+$signed( -{ 1'b0,x308 } )+$signed( -{ 1'b0,x564 } )+$signed( { 2'b0,x53 } <<<3'd1 )+$signed( -{ 1'b0,x309 } )+$signed( -{ 2'b0,x565 }<<<3'd1 )+$signed(11'd40);
assign y202=temp_y[202][11] ==1'b1 ? 5'd0 :  
        temp_y[202][8] ==1'b1 ? 5'd31 : 
        temp_y[202][2]==1'b1 ? temp_y[202][7:3]+1'b1 : temp_y[202][7:3];
assign temp_y[266] = 
+$signed( -{ 1'b0,x36 } )+$signed( { 2'b0,x292 } <<<3'd1 )+$signed( -{ 1'b0,x548 } )+$signed( -{ 1'b0,x37 } )+$signed( { 2'b0,x293 } <<<3'd1 )+$signed( -{ 2'b0,x549 }<<<3'd1 )+$signed( -{ 1'b0,x52 } )+$signed( { 2'b0,x308 } <<<3'd1 )+$signed( -{ 1'b0,x564 } )+$signed( -{ 2'b0,x53 }<<<3'd1 )+$signed( { 3'b0,x309 }<<<3'd2 )+$signed( -{ 2'b0,x565 }<<<3'd1 )+$signed(11'd32);
assign y266=temp_y[266][11] ==1'b1 ? 5'd0 :  
        temp_y[266][8] ==1'b1 ? 5'd31 : 
        temp_y[266][2]==1'b1 ? temp_y[266][7:3]+1'b1 : temp_y[266][7:3];
assign temp_y[330] = 
+$signed( -{ 1'b0,x36 } )+$signed( -{ 2'b0,x292 }<<<3'd1 )+$signed( -{ 1'b0,x548 } )+$signed( { 1'b0,x37 }  )+$signed( { 2'b0,x293 } <<<3'd1 )+$signed( { 1'b0,x549 }  )+$signed( { 1'b0,x52 }  )+$signed( { 2'b0,x308 } <<<3'd1 )+$signed( { 2'b0,x564 } <<<3'd1 )+$signed( -{ 1'b0,x53 } )+$signed( -{ 2'b0,x309 }<<<3'd1 )+$signed( -{ 1'b0,x565 } )-$signed(11'd68);
assign y330=temp_y[330][11] ==1'b1 ? 5'd0 :  
        temp_y[330][8] ==1'b1 ? 5'd31 : 
        temp_y[330][2]==1'b1 ? temp_y[330][7:3]+1'b1 : temp_y[330][7:3];
assign temp_y[394] = 
+$signed( { 1'b0,x292 }  )+$signed( { 1'b0,x549 }  )+$signed( { 1'b0,x565 }  )-$signed(11'd108);
assign y394=temp_y[394][11] ==1'b1 ? 5'd0 :  
        temp_y[394][8] ==1'b1 ? 5'd31 : 
        temp_y[394][2]==1'b1 ? temp_y[394][7:3]+1'b1 : temp_y[394][7:3];
assign temp_y[458] = 
+$signed( -{ 2'b0,x36 }<<<3'd1 )+$signed( { 2'b0,x548 } <<<3'd1 )+$signed( -{ 2'b0,x37 }<<<3'd1 )+$signed( { 1'b0,x293 }  )+$signed( { 1'b0,x549 }  )+$signed( -{ 2'b0,x52 }<<<3'd1 )+$signed( { 1'b0,x308 }  )+$signed( { 1'b0,x564 }  )+$signed( -{ 1'b0,x53 } )+$signed(11'd64);
assign y458=temp_y[458][11] ==1'b1 ? 5'd0 :  
        temp_y[458][8] ==1'b1 ? 5'd31 : 
        temp_y[458][2]==1'b1 ? temp_y[458][7:3]+1'b1 : temp_y[458][7:3];
assign temp_y[522] = 
+$signed( -{ 2'b0,x36 }<<<3'd1 )+$signed( -{ 1'b0,x292 } )+$signed( -{ 3'b0,x37 }<<<3'd2)+$signed( { 1'b0,x52 }  )+$signed( { 1'b0,x308 }  )+$signed( { 3'b0,x53 }<<<3'd2 )+$signed(11'd16);
assign y522=temp_y[522][11] ==1'b1 ? 5'd0 :  
        temp_y[522][8] ==1'b1 ? 5'd31 : 
        temp_y[522][2]==1'b1 ? temp_y[522][7:3]+1'b1 : temp_y[522][7:3];
assign temp_y[586] = 
+$signed( { 2'b0,x292 } <<<3'd1 )+$signed( { 2'b0,x548 } <<<3'd1 )+$signed( -{ 1'b0,x37 } )+$signed( -{ 2'b0,x293 }<<<3'd1 )+$signed( -{ 2'b0,x549 }<<<3'd1 )+$signed( { 2'b0,x308 } <<<3'd1 )+$signed( { 1'b0,x564 }  )+$signed( -{ 2'b0,x309 }<<<3'd1 )-$signed(11'd8);
assign y586=temp_y[586][11] ==1'b1 ? 5'd0 :  
        temp_y[586][8] ==1'b1 ? 5'd31 : 
        temp_y[586][2]==1'b1 ? temp_y[586][7:3]+1'b1 : temp_y[586][7:3];
assign temp_y[11] = 
+$signed( -{ 2'b0,x294 }<<<3'd1 )+$signed( -{ 1'b0,x550 } )+$signed( { 1'b0,x39 }  )+$signed( { 1'b0,x295 }  )+$signed( { 1'b0,x551 }  )+$signed( -{ 2'b0,x310 }<<<3'd1 )+$signed( -{ 2'b0,x566 }<<<3'd1 )+$signed( { 2'b0,x311 } <<<3'd1 )+$signed( { 2'b0,x567 } <<<3'd1 )-$signed(11'd16);
assign y11=temp_y[11][11] ==1'b1 ? 5'd0 :  
        temp_y[11][8] ==1'b1 ? 5'd31 : 
        temp_y[11][2]==1'b1 ? temp_y[11][7:3]+1'b1 : temp_y[11][7:3];
assign temp_y[75] = 
+$signed( { 3'b0,x38 }<<<3'd2 )+$signed( -{ 2'b0,x294 }<<<3'd1 )+$signed( -{ 2'b0,x550 }<<<3'd1 )+$signed( { 2'b0,x39 } <<<3'd1 )+$signed( -{ 3'b0,x295 }<<<3'd2)+$signed( { 1'b0,x551 }  )+$signed( -{ 1'b0,x54 } )+$signed( { 1'b0,x566 }  )+$signed( -{ 2'b0,x55 }<<<3'd1 )+$signed( -{ 1'b0,x311 } )+$signed( { 2'b0,x567 } <<<3'd1 )+$signed(11'd24);
assign y75=temp_y[75][11] ==1'b1 ? 5'd0 :  
        temp_y[75][8] ==1'b1 ? 5'd31 : 
        temp_y[75][2]==1'b1 ? temp_y[75][7:3]+1'b1 : temp_y[75][7:3];
assign temp_y[139] = 
+$signed( { 2'b0,x38 } <<<3'd1 )+$signed( { 2'b0,x294 } <<<3'd1 )+$signed( { 1'b0,x550 }  )+$signed( { 2'b0,x39 } <<<3'd1 )+$signed( -{ 1'b0,x295 } )+$signed( { 1'b0,x551 }  )+$signed( -{ 2'b0,x54 }<<<3'd1 )+$signed( -{ 2'b0,x310 }<<<3'd1 )+$signed( -{ 1'b0,x566 } )+$signed( -{ 1'b0,x55 } )+$signed( -{ 1'b0,x311 } )+$signed( -{ 1'b0,x567 } )+$signed(11'd16);
assign y139=temp_y[139][11] ==1'b1 ? 5'd0 :  
        temp_y[139][8] ==1'b1 ? 5'd31 : 
        temp_y[139][2]==1'b1 ? temp_y[139][7:3]+1'b1 : temp_y[139][7:3];
assign temp_y[203] = 
+$signed( { 1'b0,x38 }  )+$signed( -{ 1'b0,x294 } )+$signed( { 1'b0,x39 }  )+$signed( -{ 1'b0,x295 } )+$signed( { 2'b0,x54 } <<<3'd1 )+$signed( -{ 1'b0,x310 } )+$signed( -{ 1'b0,x566 } )+$signed( { 2'b0,x55 } <<<3'd1 )+$signed( -{ 1'b0,x311 } )+$signed( -{ 2'b0,x567 }<<<3'd1 )+$signed(11'd40);
assign y203=temp_y[203][11] ==1'b1 ? 5'd0 :  
        temp_y[203][8] ==1'b1 ? 5'd31 : 
        temp_y[203][2]==1'b1 ? temp_y[203][7:3]+1'b1 : temp_y[203][7:3];
assign temp_y[267] = 
+$signed( -{ 1'b0,x38 } )+$signed( { 2'b0,x294 } <<<3'd1 )+$signed( -{ 1'b0,x550 } )+$signed( -{ 1'b0,x39 } )+$signed( { 2'b0,x295 } <<<3'd1 )+$signed( -{ 2'b0,x551 }<<<3'd1 )+$signed( -{ 1'b0,x54 } )+$signed( { 2'b0,x310 } <<<3'd1 )+$signed( -{ 1'b0,x566 } )+$signed( -{ 2'b0,x55 }<<<3'd1 )+$signed( { 3'b0,x311 }<<<3'd2 )+$signed( -{ 2'b0,x567 }<<<3'd1 )+$signed(11'd32);
assign y267=temp_y[267][11] ==1'b1 ? 5'd0 :  
        temp_y[267][8] ==1'b1 ? 5'd31 : 
        temp_y[267][2]==1'b1 ? temp_y[267][7:3]+1'b1 : temp_y[267][7:3];
assign temp_y[331] = 
+$signed( -{ 1'b0,x38 } )+$signed( -{ 2'b0,x294 }<<<3'd1 )+$signed( -{ 1'b0,x550 } )+$signed( { 1'b0,x39 }  )+$signed( { 2'b0,x295 } <<<3'd1 )+$signed( { 1'b0,x551 }  )+$signed( { 1'b0,x54 }  )+$signed( { 2'b0,x310 } <<<3'd1 )+$signed( { 2'b0,x566 } <<<3'd1 )+$signed( -{ 1'b0,x55 } )+$signed( -{ 2'b0,x311 }<<<3'd1 )+$signed( -{ 1'b0,x567 } )-$signed(11'd68);
assign y331=temp_y[331][11] ==1'b1 ? 5'd0 :  
        temp_y[331][8] ==1'b1 ? 5'd31 : 
        temp_y[331][2]==1'b1 ? temp_y[331][7:3]+1'b1 : temp_y[331][7:3];
assign temp_y[395] = 
+$signed( { 1'b0,x294 }  )+$signed( { 1'b0,x551 }  )+$signed( { 1'b0,x567 }  )-$signed(11'd108);
assign y395=temp_y[395][11] ==1'b1 ? 5'd0 :  
        temp_y[395][8] ==1'b1 ? 5'd31 : 
        temp_y[395][2]==1'b1 ? temp_y[395][7:3]+1'b1 : temp_y[395][7:3];
assign temp_y[459] = 
+$signed( -{ 2'b0,x38 }<<<3'd1 )+$signed( { 2'b0,x550 } <<<3'd1 )+$signed( -{ 2'b0,x39 }<<<3'd1 )+$signed( { 1'b0,x295 }  )+$signed( { 1'b0,x551 }  )+$signed( -{ 2'b0,x54 }<<<3'd1 )+$signed( { 1'b0,x310 }  )+$signed( { 1'b0,x566 }  )+$signed( -{ 1'b0,x55 } )+$signed(11'd64);
assign y459=temp_y[459][11] ==1'b1 ? 5'd0 :  
        temp_y[459][8] ==1'b1 ? 5'd31 : 
        temp_y[459][2]==1'b1 ? temp_y[459][7:3]+1'b1 : temp_y[459][7:3];
assign temp_y[523] = 
+$signed( -{ 2'b0,x38 }<<<3'd1 )+$signed( -{ 1'b0,x294 } )+$signed( -{ 3'b0,x39 }<<<3'd2)+$signed( { 1'b0,x54 }  )+$signed( { 1'b0,x310 }  )+$signed( { 3'b0,x55 }<<<3'd2 )+$signed(11'd16);
assign y523=temp_y[523][11] ==1'b1 ? 5'd0 :  
        temp_y[523][8] ==1'b1 ? 5'd31 : 
        temp_y[523][2]==1'b1 ? temp_y[523][7:3]+1'b1 : temp_y[523][7:3];
assign temp_y[587] = 
+$signed( { 2'b0,x294 } <<<3'd1 )+$signed( { 2'b0,x550 } <<<3'd1 )+$signed( -{ 1'b0,x39 } )+$signed( -{ 2'b0,x295 }<<<3'd1 )+$signed( -{ 2'b0,x551 }<<<3'd1 )+$signed( { 2'b0,x310 } <<<3'd1 )+$signed( { 1'b0,x566 }  )+$signed( -{ 2'b0,x311 }<<<3'd1 )-$signed(11'd8);
assign y587=temp_y[587][11] ==1'b1 ? 5'd0 :  
        temp_y[587][8] ==1'b1 ? 5'd31 : 
        temp_y[587][2]==1'b1 ? temp_y[587][7:3]+1'b1 : temp_y[587][7:3];
assign temp_y[12] = 
+$signed( -{ 2'b0,x296 }<<<3'd1 )+$signed( -{ 1'b0,x552 } )+$signed( { 1'b0,x41 }  )+$signed( { 1'b0,x297 }  )+$signed( { 1'b0,x553 }  )+$signed( -{ 2'b0,x312 }<<<3'd1 )+$signed( -{ 2'b0,x568 }<<<3'd1 )+$signed( { 2'b0,x313 } <<<3'd1 )+$signed( { 2'b0,x569 } <<<3'd1 )-$signed(11'd16);
assign y12=temp_y[12][11] ==1'b1 ? 5'd0 :  
        temp_y[12][8] ==1'b1 ? 5'd31 : 
        temp_y[12][2]==1'b1 ? temp_y[12][7:3]+1'b1 : temp_y[12][7:3];
assign temp_y[76] = 
+$signed( { 3'b0,x40 }<<<3'd2 )+$signed( -{ 2'b0,x296 }<<<3'd1 )+$signed( -{ 2'b0,x552 }<<<3'd1 )+$signed( { 2'b0,x41 } <<<3'd1 )+$signed( -{ 3'b0,x297 }<<<3'd2)+$signed( { 1'b0,x553 }  )+$signed( -{ 1'b0,x56 } )+$signed( { 1'b0,x568 }  )+$signed( -{ 2'b0,x57 }<<<3'd1 )+$signed( -{ 1'b0,x313 } )+$signed( { 2'b0,x569 } <<<3'd1 )+$signed(11'd24);
assign y76=temp_y[76][11] ==1'b1 ? 5'd0 :  
        temp_y[76][8] ==1'b1 ? 5'd31 : 
        temp_y[76][2]==1'b1 ? temp_y[76][7:3]+1'b1 : temp_y[76][7:3];
assign temp_y[140] = 
+$signed( { 2'b0,x40 } <<<3'd1 )+$signed( { 2'b0,x296 } <<<3'd1 )+$signed( { 1'b0,x552 }  )+$signed( { 2'b0,x41 } <<<3'd1 )+$signed( -{ 1'b0,x297 } )+$signed( { 1'b0,x553 }  )+$signed( -{ 2'b0,x56 }<<<3'd1 )+$signed( -{ 2'b0,x312 }<<<3'd1 )+$signed( -{ 1'b0,x568 } )+$signed( -{ 1'b0,x57 } )+$signed( -{ 1'b0,x313 } )+$signed( -{ 1'b0,x569 } )+$signed(11'd16);
assign y140=temp_y[140][11] ==1'b1 ? 5'd0 :  
        temp_y[140][8] ==1'b1 ? 5'd31 : 
        temp_y[140][2]==1'b1 ? temp_y[140][7:3]+1'b1 : temp_y[140][7:3];
assign temp_y[204] = 
+$signed( { 1'b0,x40 }  )+$signed( -{ 1'b0,x296 } )+$signed( { 1'b0,x41 }  )+$signed( -{ 1'b0,x297 } )+$signed( { 2'b0,x56 } <<<3'd1 )+$signed( -{ 1'b0,x312 } )+$signed( -{ 1'b0,x568 } )+$signed( { 2'b0,x57 } <<<3'd1 )+$signed( -{ 1'b0,x313 } )+$signed( -{ 2'b0,x569 }<<<3'd1 )+$signed(11'd40);
assign y204=temp_y[204][11] ==1'b1 ? 5'd0 :  
        temp_y[204][8] ==1'b1 ? 5'd31 : 
        temp_y[204][2]==1'b1 ? temp_y[204][7:3]+1'b1 : temp_y[204][7:3];
assign temp_y[268] = 
+$signed( -{ 1'b0,x40 } )+$signed( { 2'b0,x296 } <<<3'd1 )+$signed( -{ 1'b0,x552 } )+$signed( -{ 1'b0,x41 } )+$signed( { 2'b0,x297 } <<<3'd1 )+$signed( -{ 2'b0,x553 }<<<3'd1 )+$signed( -{ 1'b0,x56 } )+$signed( { 2'b0,x312 } <<<3'd1 )+$signed( -{ 1'b0,x568 } )+$signed( -{ 2'b0,x57 }<<<3'd1 )+$signed( { 3'b0,x313 }<<<3'd2 )+$signed( -{ 2'b0,x569 }<<<3'd1 )+$signed(11'd32);
assign y268=temp_y[268][11] ==1'b1 ? 5'd0 :  
        temp_y[268][8] ==1'b1 ? 5'd31 : 
        temp_y[268][2]==1'b1 ? temp_y[268][7:3]+1'b1 : temp_y[268][7:3];
assign temp_y[332] = 
+$signed( -{ 1'b0,x40 } )+$signed( -{ 2'b0,x296 }<<<3'd1 )+$signed( -{ 1'b0,x552 } )+$signed( { 1'b0,x41 }  )+$signed( { 2'b0,x297 } <<<3'd1 )+$signed( { 1'b0,x553 }  )+$signed( { 1'b0,x56 }  )+$signed( { 2'b0,x312 } <<<3'd1 )+$signed( { 2'b0,x568 } <<<3'd1 )+$signed( -{ 1'b0,x57 } )+$signed( -{ 2'b0,x313 }<<<3'd1 )+$signed( -{ 1'b0,x569 } )-$signed(11'd68);
assign y332=temp_y[332][11] ==1'b1 ? 5'd0 :  
        temp_y[332][8] ==1'b1 ? 5'd31 : 
        temp_y[332][2]==1'b1 ? temp_y[332][7:3]+1'b1 : temp_y[332][7:3];
assign temp_y[396] = 
+$signed( { 1'b0,x296 }  )+$signed( { 1'b0,x553 }  )+$signed( { 1'b0,x569 }  )-$signed(11'd108);
assign y396=temp_y[396][11] ==1'b1 ? 5'd0 :  
        temp_y[396][8] ==1'b1 ? 5'd31 : 
        temp_y[396][2]==1'b1 ? temp_y[396][7:3]+1'b1 : temp_y[396][7:3];
assign temp_y[460] = 
+$signed( -{ 2'b0,x40 }<<<3'd1 )+$signed( { 2'b0,x552 } <<<3'd1 )+$signed( -{ 2'b0,x41 }<<<3'd1 )+$signed( { 1'b0,x297 }  )+$signed( { 1'b0,x553 }  )+$signed( -{ 2'b0,x56 }<<<3'd1 )+$signed( { 1'b0,x312 }  )+$signed( { 1'b0,x568 }  )+$signed( -{ 1'b0,x57 } )+$signed(11'd64);
assign y460=temp_y[460][11] ==1'b1 ? 5'd0 :  
        temp_y[460][8] ==1'b1 ? 5'd31 : 
        temp_y[460][2]==1'b1 ? temp_y[460][7:3]+1'b1 : temp_y[460][7:3];
assign temp_y[524] = 
+$signed( -{ 2'b0,x40 }<<<3'd1 )+$signed( -{ 1'b0,x296 } )+$signed( -{ 3'b0,x41 }<<<3'd2)+$signed( { 1'b0,x56 }  )+$signed( { 1'b0,x312 }  )+$signed( { 3'b0,x57 }<<<3'd2 )+$signed(11'd16);
assign y524=temp_y[524][11] ==1'b1 ? 5'd0 :  
        temp_y[524][8] ==1'b1 ? 5'd31 : 
        temp_y[524][2]==1'b1 ? temp_y[524][7:3]+1'b1 : temp_y[524][7:3];
assign temp_y[588] = 
+$signed( { 2'b0,x296 } <<<3'd1 )+$signed( { 2'b0,x552 } <<<3'd1 )+$signed( -{ 1'b0,x41 } )+$signed( -{ 2'b0,x297 }<<<3'd1 )+$signed( -{ 2'b0,x553 }<<<3'd1 )+$signed( { 2'b0,x312 } <<<3'd1 )+$signed( { 1'b0,x568 }  )+$signed( -{ 2'b0,x313 }<<<3'd1 )-$signed(11'd8);
assign y588=temp_y[588][11] ==1'b1 ? 5'd0 :  
        temp_y[588][8] ==1'b1 ? 5'd31 : 
        temp_y[588][2]==1'b1 ? temp_y[588][7:3]+1'b1 : temp_y[588][7:3];
assign temp_y[13] = 
+$signed( -{ 2'b0,x298 }<<<3'd1 )+$signed( -{ 1'b0,x554 } )+$signed( { 1'b0,x43 }  )+$signed( { 1'b0,x299 }  )+$signed( { 1'b0,x555 }  )+$signed( -{ 2'b0,x314 }<<<3'd1 )+$signed( -{ 2'b0,x570 }<<<3'd1 )+$signed( { 2'b0,x315 } <<<3'd1 )+$signed( { 2'b0,x571 } <<<3'd1 )-$signed(11'd16);
assign y13=temp_y[13][11] ==1'b1 ? 5'd0 :  
        temp_y[13][8] ==1'b1 ? 5'd31 : 
        temp_y[13][2]==1'b1 ? temp_y[13][7:3]+1'b1 : temp_y[13][7:3];
assign temp_y[77] = 
+$signed( { 3'b0,x42 }<<<3'd2 )+$signed( -{ 2'b0,x298 }<<<3'd1 )+$signed( -{ 2'b0,x554 }<<<3'd1 )+$signed( { 2'b0,x43 } <<<3'd1 )+$signed( -{ 3'b0,x299 }<<<3'd2)+$signed( { 1'b0,x555 }  )+$signed( -{ 1'b0,x58 } )+$signed( { 1'b0,x570 }  )+$signed( -{ 2'b0,x59 }<<<3'd1 )+$signed( -{ 1'b0,x315 } )+$signed( { 2'b0,x571 } <<<3'd1 )+$signed(11'd24);
assign y77=temp_y[77][11] ==1'b1 ? 5'd0 :  
        temp_y[77][8] ==1'b1 ? 5'd31 : 
        temp_y[77][2]==1'b1 ? temp_y[77][7:3]+1'b1 : temp_y[77][7:3];
assign temp_y[141] = 
+$signed( { 2'b0,x42 } <<<3'd1 )+$signed( { 2'b0,x298 } <<<3'd1 )+$signed( { 1'b0,x554 }  )+$signed( { 2'b0,x43 } <<<3'd1 )+$signed( -{ 1'b0,x299 } )+$signed( { 1'b0,x555 }  )+$signed( -{ 2'b0,x58 }<<<3'd1 )+$signed( -{ 2'b0,x314 }<<<3'd1 )+$signed( -{ 1'b0,x570 } )+$signed( -{ 1'b0,x59 } )+$signed( -{ 1'b0,x315 } )+$signed( -{ 1'b0,x571 } )+$signed(11'd16);
assign y141=temp_y[141][11] ==1'b1 ? 5'd0 :  
        temp_y[141][8] ==1'b1 ? 5'd31 : 
        temp_y[141][2]==1'b1 ? temp_y[141][7:3]+1'b1 : temp_y[141][7:3];
assign temp_y[205] = 
+$signed( { 1'b0,x42 }  )+$signed( -{ 1'b0,x298 } )+$signed( { 1'b0,x43 }  )+$signed( -{ 1'b0,x299 } )+$signed( { 2'b0,x58 } <<<3'd1 )+$signed( -{ 1'b0,x314 } )+$signed( -{ 1'b0,x570 } )+$signed( { 2'b0,x59 } <<<3'd1 )+$signed( -{ 1'b0,x315 } )+$signed( -{ 2'b0,x571 }<<<3'd1 )+$signed(11'd40);
assign y205=temp_y[205][11] ==1'b1 ? 5'd0 :  
        temp_y[205][8] ==1'b1 ? 5'd31 : 
        temp_y[205][2]==1'b1 ? temp_y[205][7:3]+1'b1 : temp_y[205][7:3];
assign temp_y[269] = 
+$signed( -{ 1'b0,x42 } )+$signed( { 2'b0,x298 } <<<3'd1 )+$signed( -{ 1'b0,x554 } )+$signed( -{ 1'b0,x43 } )+$signed( { 2'b0,x299 } <<<3'd1 )+$signed( -{ 2'b0,x555 }<<<3'd1 )+$signed( -{ 1'b0,x58 } )+$signed( { 2'b0,x314 } <<<3'd1 )+$signed( -{ 1'b0,x570 } )+$signed( -{ 2'b0,x59 }<<<3'd1 )+$signed( { 3'b0,x315 }<<<3'd2 )+$signed( -{ 2'b0,x571 }<<<3'd1 )+$signed(11'd32);
assign y269=temp_y[269][11] ==1'b1 ? 5'd0 :  
        temp_y[269][8] ==1'b1 ? 5'd31 : 
        temp_y[269][2]==1'b1 ? temp_y[269][7:3]+1'b1 : temp_y[269][7:3];
assign temp_y[333] = 
+$signed( -{ 1'b0,x42 } )+$signed( -{ 2'b0,x298 }<<<3'd1 )+$signed( -{ 1'b0,x554 } )+$signed( { 1'b0,x43 }  )+$signed( { 2'b0,x299 } <<<3'd1 )+$signed( { 1'b0,x555 }  )+$signed( { 1'b0,x58 }  )+$signed( { 2'b0,x314 } <<<3'd1 )+$signed( { 2'b0,x570 } <<<3'd1 )+$signed( -{ 1'b0,x59 } )+$signed( -{ 2'b0,x315 }<<<3'd1 )+$signed( -{ 1'b0,x571 } )-$signed(11'd68);
assign y333=temp_y[333][11] ==1'b1 ? 5'd0 :  
        temp_y[333][8] ==1'b1 ? 5'd31 : 
        temp_y[333][2]==1'b1 ? temp_y[333][7:3]+1'b1 : temp_y[333][7:3];
assign temp_y[397] = 
+$signed( { 1'b0,x298 }  )+$signed( { 1'b0,x555 }  )+$signed( { 1'b0,x571 }  )-$signed(11'd108);
assign y397=temp_y[397][11] ==1'b1 ? 5'd0 :  
        temp_y[397][8] ==1'b1 ? 5'd31 : 
        temp_y[397][2]==1'b1 ? temp_y[397][7:3]+1'b1 : temp_y[397][7:3];
assign temp_y[461] = 
+$signed( -{ 2'b0,x42 }<<<3'd1 )+$signed( { 2'b0,x554 } <<<3'd1 )+$signed( -{ 2'b0,x43 }<<<3'd1 )+$signed( { 1'b0,x299 }  )+$signed( { 1'b0,x555 }  )+$signed( -{ 2'b0,x58 }<<<3'd1 )+$signed( { 1'b0,x314 }  )+$signed( { 1'b0,x570 }  )+$signed( -{ 1'b0,x59 } )+$signed(11'd64);
assign y461=temp_y[461][11] ==1'b1 ? 5'd0 :  
        temp_y[461][8] ==1'b1 ? 5'd31 : 
        temp_y[461][2]==1'b1 ? temp_y[461][7:3]+1'b1 : temp_y[461][7:3];
assign temp_y[525] = 
+$signed( -{ 2'b0,x42 }<<<3'd1 )+$signed( -{ 1'b0,x298 } )+$signed( -{ 3'b0,x43 }<<<3'd2)+$signed( { 1'b0,x58 }  )+$signed( { 1'b0,x314 }  )+$signed( { 3'b0,x59 }<<<3'd2 )+$signed(11'd16);
assign y525=temp_y[525][11] ==1'b1 ? 5'd0 :  
        temp_y[525][8] ==1'b1 ? 5'd31 : 
        temp_y[525][2]==1'b1 ? temp_y[525][7:3]+1'b1 : temp_y[525][7:3];
assign temp_y[589] = 
+$signed( { 2'b0,x298 } <<<3'd1 )+$signed( { 2'b0,x554 } <<<3'd1 )+$signed( -{ 1'b0,x43 } )+$signed( -{ 2'b0,x299 }<<<3'd1 )+$signed( -{ 2'b0,x555 }<<<3'd1 )+$signed( { 2'b0,x314 } <<<3'd1 )+$signed( { 1'b0,x570 }  )+$signed( -{ 2'b0,x315 }<<<3'd1 )-$signed(11'd8);
assign y589=temp_y[589][11] ==1'b1 ? 5'd0 :  
        temp_y[589][8] ==1'b1 ? 5'd31 : 
        temp_y[589][2]==1'b1 ? temp_y[589][7:3]+1'b1 : temp_y[589][7:3];
assign temp_y[14] = 
+$signed( -{ 2'b0,x300 }<<<3'd1 )+$signed( -{ 1'b0,x556 } )+$signed( { 1'b0,x45 }  )+$signed( { 1'b0,x301 }  )+$signed( { 1'b0,x557 }  )+$signed( -{ 2'b0,x316 }<<<3'd1 )+$signed( -{ 2'b0,x572 }<<<3'd1 )+$signed( { 2'b0,x317 } <<<3'd1 )+$signed( { 2'b0,x573 } <<<3'd1 )-$signed(11'd16);
assign y14=temp_y[14][11] ==1'b1 ? 5'd0 :  
        temp_y[14][8] ==1'b1 ? 5'd31 : 
        temp_y[14][2]==1'b1 ? temp_y[14][7:3]+1'b1 : temp_y[14][7:3];
assign temp_y[78] = 
+$signed( { 3'b0,x44 }<<<3'd2 )+$signed( -{ 2'b0,x300 }<<<3'd1 )+$signed( -{ 2'b0,x556 }<<<3'd1 )+$signed( { 2'b0,x45 } <<<3'd1 )+$signed( -{ 3'b0,x301 }<<<3'd2)+$signed( { 1'b0,x557 }  )+$signed( -{ 1'b0,x60 } )+$signed( { 1'b0,x572 }  )+$signed( -{ 2'b0,x61 }<<<3'd1 )+$signed( -{ 1'b0,x317 } )+$signed( { 2'b0,x573 } <<<3'd1 )+$signed(11'd24);
assign y78=temp_y[78][11] ==1'b1 ? 5'd0 :  
        temp_y[78][8] ==1'b1 ? 5'd31 : 
        temp_y[78][2]==1'b1 ? temp_y[78][7:3]+1'b1 : temp_y[78][7:3];
assign temp_y[142] = 
+$signed( { 2'b0,x44 } <<<3'd1 )+$signed( { 2'b0,x300 } <<<3'd1 )+$signed( { 1'b0,x556 }  )+$signed( { 2'b0,x45 } <<<3'd1 )+$signed( -{ 1'b0,x301 } )+$signed( { 1'b0,x557 }  )+$signed( -{ 2'b0,x60 }<<<3'd1 )+$signed( -{ 2'b0,x316 }<<<3'd1 )+$signed( -{ 1'b0,x572 } )+$signed( -{ 1'b0,x61 } )+$signed( -{ 1'b0,x317 } )+$signed( -{ 1'b0,x573 } )+$signed(11'd16);
assign y142=temp_y[142][11] ==1'b1 ? 5'd0 :  
        temp_y[142][8] ==1'b1 ? 5'd31 : 
        temp_y[142][2]==1'b1 ? temp_y[142][7:3]+1'b1 : temp_y[142][7:3];
assign temp_y[206] = 
+$signed( { 1'b0,x44 }  )+$signed( -{ 1'b0,x300 } )+$signed( { 1'b0,x45 }  )+$signed( -{ 1'b0,x301 } )+$signed( { 2'b0,x60 } <<<3'd1 )+$signed( -{ 1'b0,x316 } )+$signed( -{ 1'b0,x572 } )+$signed( { 2'b0,x61 } <<<3'd1 )+$signed( -{ 1'b0,x317 } )+$signed( -{ 2'b0,x573 }<<<3'd1 )+$signed(11'd40);
assign y206=temp_y[206][11] ==1'b1 ? 5'd0 :  
        temp_y[206][8] ==1'b1 ? 5'd31 : 
        temp_y[206][2]==1'b1 ? temp_y[206][7:3]+1'b1 : temp_y[206][7:3];
assign temp_y[270] = 
+$signed( -{ 1'b0,x44 } )+$signed( { 2'b0,x300 } <<<3'd1 )+$signed( -{ 1'b0,x556 } )+$signed( -{ 1'b0,x45 } )+$signed( { 2'b0,x301 } <<<3'd1 )+$signed( -{ 2'b0,x557 }<<<3'd1 )+$signed( -{ 1'b0,x60 } )+$signed( { 2'b0,x316 } <<<3'd1 )+$signed( -{ 1'b0,x572 } )+$signed( -{ 2'b0,x61 }<<<3'd1 )+$signed( { 3'b0,x317 }<<<3'd2 )+$signed( -{ 2'b0,x573 }<<<3'd1 )+$signed(11'd32);
assign y270=temp_y[270][11] ==1'b1 ? 5'd0 :  
        temp_y[270][8] ==1'b1 ? 5'd31 : 
        temp_y[270][2]==1'b1 ? temp_y[270][7:3]+1'b1 : temp_y[270][7:3];
assign temp_y[334] = 
+$signed( -{ 1'b0,x44 } )+$signed( -{ 2'b0,x300 }<<<3'd1 )+$signed( -{ 1'b0,x556 } )+$signed( { 1'b0,x45 }  )+$signed( { 2'b0,x301 } <<<3'd1 )+$signed( { 1'b0,x557 }  )+$signed( { 1'b0,x60 }  )+$signed( { 2'b0,x316 } <<<3'd1 )+$signed( { 2'b0,x572 } <<<3'd1 )+$signed( -{ 1'b0,x61 } )+$signed( -{ 2'b0,x317 }<<<3'd1 )+$signed( -{ 1'b0,x573 } )-$signed(11'd68);
assign y334=temp_y[334][11] ==1'b1 ? 5'd0 :  
        temp_y[334][8] ==1'b1 ? 5'd31 : 
        temp_y[334][2]==1'b1 ? temp_y[334][7:3]+1'b1 : temp_y[334][7:3];
assign temp_y[398] = 
+$signed( { 1'b0,x300 }  )+$signed( { 1'b0,x557 }  )+$signed( { 1'b0,x573 }  )-$signed(11'd108);
assign y398=temp_y[398][11] ==1'b1 ? 5'd0 :  
        temp_y[398][8] ==1'b1 ? 5'd31 : 
        temp_y[398][2]==1'b1 ? temp_y[398][7:3]+1'b1 : temp_y[398][7:3];
assign temp_y[462] = 
+$signed( -{ 2'b0,x44 }<<<3'd1 )+$signed( { 2'b0,x556 } <<<3'd1 )+$signed( -{ 2'b0,x45 }<<<3'd1 )+$signed( { 1'b0,x301 }  )+$signed( { 1'b0,x557 }  )+$signed( -{ 2'b0,x60 }<<<3'd1 )+$signed( { 1'b0,x316 }  )+$signed( { 1'b0,x572 }  )+$signed( -{ 1'b0,x61 } )+$signed(11'd64);
assign y462=temp_y[462][11] ==1'b1 ? 5'd0 :  
        temp_y[462][8] ==1'b1 ? 5'd31 : 
        temp_y[462][2]==1'b1 ? temp_y[462][7:3]+1'b1 : temp_y[462][7:3];
assign temp_y[526] = 
+$signed( -{ 2'b0,x44 }<<<3'd1 )+$signed( -{ 1'b0,x300 } )+$signed( -{ 3'b0,x45 }<<<3'd2)+$signed( { 1'b0,x60 }  )+$signed( { 1'b0,x316 }  )+$signed( { 3'b0,x61 }<<<3'd2 )+$signed(11'd16);
assign y526=temp_y[526][11] ==1'b1 ? 5'd0 :  
        temp_y[526][8] ==1'b1 ? 5'd31 : 
        temp_y[526][2]==1'b1 ? temp_y[526][7:3]+1'b1 : temp_y[526][7:3];
assign temp_y[590] = 
+$signed( { 2'b0,x300 } <<<3'd1 )+$signed( { 2'b0,x556 } <<<3'd1 )+$signed( -{ 1'b0,x45 } )+$signed( -{ 2'b0,x301 }<<<3'd1 )+$signed( -{ 2'b0,x557 }<<<3'd1 )+$signed( { 2'b0,x316 } <<<3'd1 )+$signed( { 1'b0,x572 }  )+$signed( -{ 2'b0,x317 }<<<3'd1 )-$signed(11'd8);
assign y590=temp_y[590][11] ==1'b1 ? 5'd0 :  
        temp_y[590][8] ==1'b1 ? 5'd31 : 
        temp_y[590][2]==1'b1 ? temp_y[590][7:3]+1'b1 : temp_y[590][7:3];
assign temp_y[15] = 
+$signed( -{ 2'b0,x302 }<<<3'd1 )+$signed( -{ 1'b0,x558 } )+$signed( { 1'b0,x47 }  )+$signed( { 1'b0,x303 }  )+$signed( { 1'b0,x559 }  )+$signed( -{ 2'b0,x318 }<<<3'd1 )+$signed( -{ 2'b0,x574 }<<<3'd1 )+$signed( { 2'b0,x319 } <<<3'd1 )+$signed( { 2'b0,x575 } <<<3'd1 )-$signed(11'd16);
assign y15=temp_y[15][11] ==1'b1 ? 5'd0 :  
        temp_y[15][8] ==1'b1 ? 5'd31 : 
        temp_y[15][2]==1'b1 ? temp_y[15][7:3]+1'b1 : temp_y[15][7:3];
assign temp_y[79] = 
+$signed( { 3'b0,x46 }<<<3'd2 )+$signed( -{ 2'b0,x302 }<<<3'd1 )+$signed( -{ 2'b0,x558 }<<<3'd1 )+$signed( { 2'b0,x47 } <<<3'd1 )+$signed( -{ 3'b0,x303 }<<<3'd2)+$signed( { 1'b0,x559 }  )+$signed( -{ 1'b0,x62 } )+$signed( { 1'b0,x574 }  )+$signed( -{ 2'b0,x63 }<<<3'd1 )+$signed( -{ 1'b0,x319 } )+$signed( { 2'b0,x575 } <<<3'd1 )+$signed(11'd24);
assign y79=temp_y[79][11] ==1'b1 ? 5'd0 :  
        temp_y[79][8] ==1'b1 ? 5'd31 : 
        temp_y[79][2]==1'b1 ? temp_y[79][7:3]+1'b1 : temp_y[79][7:3];
assign temp_y[143] = 
+$signed( { 2'b0,x46 } <<<3'd1 )+$signed( { 2'b0,x302 } <<<3'd1 )+$signed( { 1'b0,x558 }  )+$signed( { 2'b0,x47 } <<<3'd1 )+$signed( -{ 1'b0,x303 } )+$signed( { 1'b0,x559 }  )+$signed( -{ 2'b0,x62 }<<<3'd1 )+$signed( -{ 2'b0,x318 }<<<3'd1 )+$signed( -{ 1'b0,x574 } )+$signed( -{ 1'b0,x63 } )+$signed( -{ 1'b0,x319 } )+$signed( -{ 1'b0,x575 } )+$signed(11'd16);
assign y143=temp_y[143][11] ==1'b1 ? 5'd0 :  
        temp_y[143][8] ==1'b1 ? 5'd31 : 
        temp_y[143][2]==1'b1 ? temp_y[143][7:3]+1'b1 : temp_y[143][7:3];
assign temp_y[207] = 
+$signed( { 1'b0,x46 }  )+$signed( -{ 1'b0,x302 } )+$signed( { 1'b0,x47 }  )+$signed( -{ 1'b0,x303 } )+$signed( { 2'b0,x62 } <<<3'd1 )+$signed( -{ 1'b0,x318 } )+$signed( -{ 1'b0,x574 } )+$signed( { 2'b0,x63 } <<<3'd1 )+$signed( -{ 1'b0,x319 } )+$signed( -{ 2'b0,x575 }<<<3'd1 )+$signed(11'd40);
assign y207=temp_y[207][11] ==1'b1 ? 5'd0 :  
        temp_y[207][8] ==1'b1 ? 5'd31 : 
        temp_y[207][2]==1'b1 ? temp_y[207][7:3]+1'b1 : temp_y[207][7:3];
assign temp_y[271] = 
+$signed( -{ 1'b0,x46 } )+$signed( { 2'b0,x302 } <<<3'd1 )+$signed( -{ 1'b0,x558 } )+$signed( -{ 1'b0,x47 } )+$signed( { 2'b0,x303 } <<<3'd1 )+$signed( -{ 2'b0,x559 }<<<3'd1 )+$signed( -{ 1'b0,x62 } )+$signed( { 2'b0,x318 } <<<3'd1 )+$signed( -{ 1'b0,x574 } )+$signed( -{ 2'b0,x63 }<<<3'd1 )+$signed( { 3'b0,x319 }<<<3'd2 )+$signed( -{ 2'b0,x575 }<<<3'd1 )+$signed(11'd32);
assign y271=temp_y[271][11] ==1'b1 ? 5'd0 :  
        temp_y[271][8] ==1'b1 ? 5'd31 : 
        temp_y[271][2]==1'b1 ? temp_y[271][7:3]+1'b1 : temp_y[271][7:3];
assign temp_y[335] = 
+$signed( -{ 1'b0,x46 } )+$signed( -{ 2'b0,x302 }<<<3'd1 )+$signed( -{ 1'b0,x558 } )+$signed( { 1'b0,x47 }  )+$signed( { 2'b0,x303 } <<<3'd1 )+$signed( { 1'b0,x559 }  )+$signed( { 1'b0,x62 }  )+$signed( { 2'b0,x318 } <<<3'd1 )+$signed( { 2'b0,x574 } <<<3'd1 )+$signed( -{ 1'b0,x63 } )+$signed( -{ 2'b0,x319 }<<<3'd1 )+$signed( -{ 1'b0,x575 } )-$signed(11'd68);
assign y335=temp_y[335][11] ==1'b1 ? 5'd0 :  
        temp_y[335][8] ==1'b1 ? 5'd31 : 
        temp_y[335][2]==1'b1 ? temp_y[335][7:3]+1'b1 : temp_y[335][7:3];
assign temp_y[399] = 
+$signed( { 1'b0,x302 }  )+$signed( { 1'b0,x559 }  )+$signed( { 1'b0,x575 }  )-$signed(11'd108);
assign y399=temp_y[399][11] ==1'b1 ? 5'd0 :  
        temp_y[399][8] ==1'b1 ? 5'd31 : 
        temp_y[399][2]==1'b1 ? temp_y[399][7:3]+1'b1 : temp_y[399][7:3];
assign temp_y[463] = 
+$signed( -{ 2'b0,x46 }<<<3'd1 )+$signed( { 2'b0,x558 } <<<3'd1 )+$signed( -{ 2'b0,x47 }<<<3'd1 )+$signed( { 1'b0,x303 }  )+$signed( { 1'b0,x559 }  )+$signed( -{ 2'b0,x62 }<<<3'd1 )+$signed( { 1'b0,x318 }  )+$signed( { 1'b0,x574 }  )+$signed( -{ 1'b0,x63 } )+$signed(11'd64);
assign y463=temp_y[463][11] ==1'b1 ? 5'd0 :  
        temp_y[463][8] ==1'b1 ? 5'd31 : 
        temp_y[463][2]==1'b1 ? temp_y[463][7:3]+1'b1 : temp_y[463][7:3];
assign temp_y[527] = 
+$signed( -{ 2'b0,x46 }<<<3'd1 )+$signed( -{ 1'b0,x302 } )+$signed( -{ 3'b0,x47 }<<<3'd2)+$signed( { 1'b0,x62 }  )+$signed( { 1'b0,x318 }  )+$signed( { 3'b0,x63 }<<<3'd2 )+$signed(11'd16);
assign y527=temp_y[527][11] ==1'b1 ? 5'd0 :  
        temp_y[527][8] ==1'b1 ? 5'd31 : 
        temp_y[527][2]==1'b1 ? temp_y[527][7:3]+1'b1 : temp_y[527][7:3];
assign temp_y[591] = 
+$signed( { 2'b0,x302 } <<<3'd1 )+$signed( { 2'b0,x558 } <<<3'd1 )+$signed( -{ 1'b0,x47 } )+$signed( -{ 2'b0,x303 }<<<3'd1 )+$signed( -{ 2'b0,x559 }<<<3'd1 )+$signed( { 2'b0,x318 } <<<3'd1 )+$signed( { 1'b0,x574 }  )+$signed( -{ 2'b0,x319 }<<<3'd1 )-$signed(11'd8);
assign y591=temp_y[591][11] ==1'b1 ? 5'd0 :  
        temp_y[591][8] ==1'b1 ? 5'd31 : 
        temp_y[591][2]==1'b1 ? temp_y[591][7:3]+1'b1 : temp_y[591][7:3];
assign temp_y[16] = 
+$signed( -{ 2'b0,x320 }<<<3'd1 )+$signed( -{ 1'b0,x576 } )+$signed( { 1'b0,x65 }  )+$signed( { 1'b0,x321 }  )+$signed( { 1'b0,x577 }  )+$signed( -{ 2'b0,x336 }<<<3'd1 )+$signed( -{ 2'b0,x592 }<<<3'd1 )+$signed( { 2'b0,x337 } <<<3'd1 )+$signed( { 2'b0,x593 } <<<3'd1 )-$signed(11'd16);
assign y16=temp_y[16][11] ==1'b1 ? 5'd0 :  
        temp_y[16][8] ==1'b1 ? 5'd31 : 
        temp_y[16][2]==1'b1 ? temp_y[16][7:3]+1'b1 : temp_y[16][7:3];
assign temp_y[80] = 
+$signed( { 3'b0,x64 }<<<3'd2 )+$signed( -{ 2'b0,x320 }<<<3'd1 )+$signed( -{ 2'b0,x576 }<<<3'd1 )+$signed( { 2'b0,x65 } <<<3'd1 )+$signed( -{ 3'b0,x321 }<<<3'd2)+$signed( { 1'b0,x577 }  )+$signed( -{ 1'b0,x80 } )+$signed( { 1'b0,x592 }  )+$signed( -{ 2'b0,x81 }<<<3'd1 )+$signed( -{ 1'b0,x337 } )+$signed( { 2'b0,x593 } <<<3'd1 )+$signed(11'd24);
assign y80=temp_y[80][11] ==1'b1 ? 5'd0 :  
        temp_y[80][8] ==1'b1 ? 5'd31 : 
        temp_y[80][2]==1'b1 ? temp_y[80][7:3]+1'b1 : temp_y[80][7:3];
assign temp_y[144] = 
+$signed( { 2'b0,x64 } <<<3'd1 )+$signed( { 2'b0,x320 } <<<3'd1 )+$signed( { 1'b0,x576 }  )+$signed( { 2'b0,x65 } <<<3'd1 )+$signed( -{ 1'b0,x321 } )+$signed( { 1'b0,x577 }  )+$signed( -{ 2'b0,x80 }<<<3'd1 )+$signed( -{ 2'b0,x336 }<<<3'd1 )+$signed( -{ 1'b0,x592 } )+$signed( -{ 1'b0,x81 } )+$signed( -{ 1'b0,x337 } )+$signed( -{ 1'b0,x593 } )+$signed(11'd16);
assign y144=temp_y[144][11] ==1'b1 ? 5'd0 :  
        temp_y[144][8] ==1'b1 ? 5'd31 : 
        temp_y[144][2]==1'b1 ? temp_y[144][7:3]+1'b1 : temp_y[144][7:3];
assign temp_y[208] = 
+$signed( { 1'b0,x64 }  )+$signed( -{ 1'b0,x320 } )+$signed( { 1'b0,x65 }  )+$signed( -{ 1'b0,x321 } )+$signed( { 2'b0,x80 } <<<3'd1 )+$signed( -{ 1'b0,x336 } )+$signed( -{ 1'b0,x592 } )+$signed( { 2'b0,x81 } <<<3'd1 )+$signed( -{ 1'b0,x337 } )+$signed( -{ 2'b0,x593 }<<<3'd1 )+$signed(11'd40);
assign y208=temp_y[208][11] ==1'b1 ? 5'd0 :  
        temp_y[208][8] ==1'b1 ? 5'd31 : 
        temp_y[208][2]==1'b1 ? temp_y[208][7:3]+1'b1 : temp_y[208][7:3];
assign temp_y[272] = 
+$signed( -{ 1'b0,x64 } )+$signed( { 2'b0,x320 } <<<3'd1 )+$signed( -{ 1'b0,x576 } )+$signed( -{ 1'b0,x65 } )+$signed( { 2'b0,x321 } <<<3'd1 )+$signed( -{ 2'b0,x577 }<<<3'd1 )+$signed( -{ 1'b0,x80 } )+$signed( { 2'b0,x336 } <<<3'd1 )+$signed( -{ 1'b0,x592 } )+$signed( -{ 2'b0,x81 }<<<3'd1 )+$signed( { 3'b0,x337 }<<<3'd2 )+$signed( -{ 2'b0,x593 }<<<3'd1 )+$signed(11'd32);
assign y272=temp_y[272][11] ==1'b1 ? 5'd0 :  
        temp_y[272][8] ==1'b1 ? 5'd31 : 
        temp_y[272][2]==1'b1 ? temp_y[272][7:3]+1'b1 : temp_y[272][7:3];
assign temp_y[336] = 
+$signed( -{ 1'b0,x64 } )+$signed( -{ 2'b0,x320 }<<<3'd1 )+$signed( -{ 1'b0,x576 } )+$signed( { 1'b0,x65 }  )+$signed( { 2'b0,x321 } <<<3'd1 )+$signed( { 1'b0,x577 }  )+$signed( { 1'b0,x80 }  )+$signed( { 2'b0,x336 } <<<3'd1 )+$signed( { 2'b0,x592 } <<<3'd1 )+$signed( -{ 1'b0,x81 } )+$signed( -{ 2'b0,x337 }<<<3'd1 )+$signed( -{ 1'b0,x593 } )-$signed(11'd68);
assign y336=temp_y[336][11] ==1'b1 ? 5'd0 :  
        temp_y[336][8] ==1'b1 ? 5'd31 : 
        temp_y[336][2]==1'b1 ? temp_y[336][7:3]+1'b1 : temp_y[336][7:3];
assign temp_y[400] = 
+$signed( { 1'b0,x320 }  )+$signed( { 1'b0,x577 }  )+$signed( { 1'b0,x593 }  )-$signed(11'd108);
assign y400=temp_y[400][11] ==1'b1 ? 5'd0 :  
        temp_y[400][8] ==1'b1 ? 5'd31 : 
        temp_y[400][2]==1'b1 ? temp_y[400][7:3]+1'b1 : temp_y[400][7:3];
assign temp_y[464] = 
+$signed( -{ 2'b0,x64 }<<<3'd1 )+$signed( { 2'b0,x576 } <<<3'd1 )+$signed( -{ 2'b0,x65 }<<<3'd1 )+$signed( { 1'b0,x321 }  )+$signed( { 1'b0,x577 }  )+$signed( -{ 2'b0,x80 }<<<3'd1 )+$signed( { 1'b0,x336 }  )+$signed( { 1'b0,x592 }  )+$signed( -{ 1'b0,x81 } )+$signed(11'd64);
assign y464=temp_y[464][11] ==1'b1 ? 5'd0 :  
        temp_y[464][8] ==1'b1 ? 5'd31 : 
        temp_y[464][2]==1'b1 ? temp_y[464][7:3]+1'b1 : temp_y[464][7:3];
assign temp_y[528] = 
+$signed( -{ 2'b0,x64 }<<<3'd1 )+$signed( -{ 1'b0,x320 } )+$signed( -{ 3'b0,x65 }<<<3'd2)+$signed( { 1'b0,x80 }  )+$signed( { 1'b0,x336 }  )+$signed( { 3'b0,x81 }<<<3'd2 )+$signed(11'd16);
assign y528=temp_y[528][11] ==1'b1 ? 5'd0 :  
        temp_y[528][8] ==1'b1 ? 5'd31 : 
        temp_y[528][2]==1'b1 ? temp_y[528][7:3]+1'b1 : temp_y[528][7:3];
assign temp_y[592] = 
+$signed( { 2'b0,x320 } <<<3'd1 )+$signed( { 2'b0,x576 } <<<3'd1 )+$signed( -{ 1'b0,x65 } )+$signed( -{ 2'b0,x321 }<<<3'd1 )+$signed( -{ 2'b0,x577 }<<<3'd1 )+$signed( { 2'b0,x336 } <<<3'd1 )+$signed( { 1'b0,x592 }  )+$signed( -{ 2'b0,x337 }<<<3'd1 )-$signed(11'd8);
assign y592=temp_y[592][11] ==1'b1 ? 5'd0 :  
        temp_y[592][8] ==1'b1 ? 5'd31 : 
        temp_y[592][2]==1'b1 ? temp_y[592][7:3]+1'b1 : temp_y[592][7:3];
assign temp_y[17] = 
+$signed( -{ 2'b0,x322 }<<<3'd1 )+$signed( -{ 1'b0,x578 } )+$signed( { 1'b0,x67 }  )+$signed( { 1'b0,x323 }  )+$signed( { 1'b0,x579 }  )+$signed( -{ 2'b0,x338 }<<<3'd1 )+$signed( -{ 2'b0,x594 }<<<3'd1 )+$signed( { 2'b0,x339 } <<<3'd1 )+$signed( { 2'b0,x595 } <<<3'd1 )-$signed(11'd16);
assign y17=temp_y[17][11] ==1'b1 ? 5'd0 :  
        temp_y[17][8] ==1'b1 ? 5'd31 : 
        temp_y[17][2]==1'b1 ? temp_y[17][7:3]+1'b1 : temp_y[17][7:3];
assign temp_y[81] = 
+$signed( { 3'b0,x66 }<<<3'd2 )+$signed( -{ 2'b0,x322 }<<<3'd1 )+$signed( -{ 2'b0,x578 }<<<3'd1 )+$signed( { 2'b0,x67 } <<<3'd1 )+$signed( -{ 3'b0,x323 }<<<3'd2)+$signed( { 1'b0,x579 }  )+$signed( -{ 1'b0,x82 } )+$signed( { 1'b0,x594 }  )+$signed( -{ 2'b0,x83 }<<<3'd1 )+$signed( -{ 1'b0,x339 } )+$signed( { 2'b0,x595 } <<<3'd1 )+$signed(11'd24);
assign y81=temp_y[81][11] ==1'b1 ? 5'd0 :  
        temp_y[81][8] ==1'b1 ? 5'd31 : 
        temp_y[81][2]==1'b1 ? temp_y[81][7:3]+1'b1 : temp_y[81][7:3];
assign temp_y[145] = 
+$signed( { 2'b0,x66 } <<<3'd1 )+$signed( { 2'b0,x322 } <<<3'd1 )+$signed( { 1'b0,x578 }  )+$signed( { 2'b0,x67 } <<<3'd1 )+$signed( -{ 1'b0,x323 } )+$signed( { 1'b0,x579 }  )+$signed( -{ 2'b0,x82 }<<<3'd1 )+$signed( -{ 2'b0,x338 }<<<3'd1 )+$signed( -{ 1'b0,x594 } )+$signed( -{ 1'b0,x83 } )+$signed( -{ 1'b0,x339 } )+$signed( -{ 1'b0,x595 } )+$signed(11'd16);
assign y145=temp_y[145][11] ==1'b1 ? 5'd0 :  
        temp_y[145][8] ==1'b1 ? 5'd31 : 
        temp_y[145][2]==1'b1 ? temp_y[145][7:3]+1'b1 : temp_y[145][7:3];
assign temp_y[209] = 
+$signed( { 1'b0,x66 }  )+$signed( -{ 1'b0,x322 } )+$signed( { 1'b0,x67 }  )+$signed( -{ 1'b0,x323 } )+$signed( { 2'b0,x82 } <<<3'd1 )+$signed( -{ 1'b0,x338 } )+$signed( -{ 1'b0,x594 } )+$signed( { 2'b0,x83 } <<<3'd1 )+$signed( -{ 1'b0,x339 } )+$signed( -{ 2'b0,x595 }<<<3'd1 )+$signed(11'd40);
assign y209=temp_y[209][11] ==1'b1 ? 5'd0 :  
        temp_y[209][8] ==1'b1 ? 5'd31 : 
        temp_y[209][2]==1'b1 ? temp_y[209][7:3]+1'b1 : temp_y[209][7:3];
assign temp_y[273] = 
+$signed( -{ 1'b0,x66 } )+$signed( { 2'b0,x322 } <<<3'd1 )+$signed( -{ 1'b0,x578 } )+$signed( -{ 1'b0,x67 } )+$signed( { 2'b0,x323 } <<<3'd1 )+$signed( -{ 2'b0,x579 }<<<3'd1 )+$signed( -{ 1'b0,x82 } )+$signed( { 2'b0,x338 } <<<3'd1 )+$signed( -{ 1'b0,x594 } )+$signed( -{ 2'b0,x83 }<<<3'd1 )+$signed( { 3'b0,x339 }<<<3'd2 )+$signed( -{ 2'b0,x595 }<<<3'd1 )+$signed(11'd32);
assign y273=temp_y[273][11] ==1'b1 ? 5'd0 :  
        temp_y[273][8] ==1'b1 ? 5'd31 : 
        temp_y[273][2]==1'b1 ? temp_y[273][7:3]+1'b1 : temp_y[273][7:3];
assign temp_y[337] = 
+$signed( -{ 1'b0,x66 } )+$signed( -{ 2'b0,x322 }<<<3'd1 )+$signed( -{ 1'b0,x578 } )+$signed( { 1'b0,x67 }  )+$signed( { 2'b0,x323 } <<<3'd1 )+$signed( { 1'b0,x579 }  )+$signed( { 1'b0,x82 }  )+$signed( { 2'b0,x338 } <<<3'd1 )+$signed( { 2'b0,x594 } <<<3'd1 )+$signed( -{ 1'b0,x83 } )+$signed( -{ 2'b0,x339 }<<<3'd1 )+$signed( -{ 1'b0,x595 } )-$signed(11'd68);
assign y337=temp_y[337][11] ==1'b1 ? 5'd0 :  
        temp_y[337][8] ==1'b1 ? 5'd31 : 
        temp_y[337][2]==1'b1 ? temp_y[337][7:3]+1'b1 : temp_y[337][7:3];
assign temp_y[401] = 
+$signed( { 1'b0,x322 }  )+$signed( { 1'b0,x579 }  )+$signed( { 1'b0,x595 }  )-$signed(11'd108);
assign y401=temp_y[401][11] ==1'b1 ? 5'd0 :  
        temp_y[401][8] ==1'b1 ? 5'd31 : 
        temp_y[401][2]==1'b1 ? temp_y[401][7:3]+1'b1 : temp_y[401][7:3];
assign temp_y[465] = 
+$signed( -{ 2'b0,x66 }<<<3'd1 )+$signed( { 2'b0,x578 } <<<3'd1 )+$signed( -{ 2'b0,x67 }<<<3'd1 )+$signed( { 1'b0,x323 }  )+$signed( { 1'b0,x579 }  )+$signed( -{ 2'b0,x82 }<<<3'd1 )+$signed( { 1'b0,x338 }  )+$signed( { 1'b0,x594 }  )+$signed( -{ 1'b0,x83 } )+$signed(11'd64);
assign y465=temp_y[465][11] ==1'b1 ? 5'd0 :  
        temp_y[465][8] ==1'b1 ? 5'd31 : 
        temp_y[465][2]==1'b1 ? temp_y[465][7:3]+1'b1 : temp_y[465][7:3];
assign temp_y[529] = 
+$signed( -{ 2'b0,x66 }<<<3'd1 )+$signed( -{ 1'b0,x322 } )+$signed( -{ 3'b0,x67 }<<<3'd2)+$signed( { 1'b0,x82 }  )+$signed( { 1'b0,x338 }  )+$signed( { 3'b0,x83 }<<<3'd2 )+$signed(11'd16);
assign y529=temp_y[529][11] ==1'b1 ? 5'd0 :  
        temp_y[529][8] ==1'b1 ? 5'd31 : 
        temp_y[529][2]==1'b1 ? temp_y[529][7:3]+1'b1 : temp_y[529][7:3];
assign temp_y[593] = 
+$signed( { 2'b0,x322 } <<<3'd1 )+$signed( { 2'b0,x578 } <<<3'd1 )+$signed( -{ 1'b0,x67 } )+$signed( -{ 2'b0,x323 }<<<3'd1 )+$signed( -{ 2'b0,x579 }<<<3'd1 )+$signed( { 2'b0,x338 } <<<3'd1 )+$signed( { 1'b0,x594 }  )+$signed( -{ 2'b0,x339 }<<<3'd1 )-$signed(11'd8);
assign y593=temp_y[593][11] ==1'b1 ? 5'd0 :  
        temp_y[593][8] ==1'b1 ? 5'd31 : 
        temp_y[593][2]==1'b1 ? temp_y[593][7:3]+1'b1 : temp_y[593][7:3];
assign temp_y[18] = 
+$signed( -{ 2'b0,x324 }<<<3'd1 )+$signed( -{ 1'b0,x580 } )+$signed( { 1'b0,x69 }  )+$signed( { 1'b0,x325 }  )+$signed( { 1'b0,x581 }  )+$signed( -{ 2'b0,x340 }<<<3'd1 )+$signed( -{ 2'b0,x596 }<<<3'd1 )+$signed( { 2'b0,x341 } <<<3'd1 )+$signed( { 2'b0,x597 } <<<3'd1 )-$signed(11'd16);
assign y18=temp_y[18][11] ==1'b1 ? 5'd0 :  
        temp_y[18][8] ==1'b1 ? 5'd31 : 
        temp_y[18][2]==1'b1 ? temp_y[18][7:3]+1'b1 : temp_y[18][7:3];
assign temp_y[82] = 
+$signed( { 3'b0,x68 }<<<3'd2 )+$signed( -{ 2'b0,x324 }<<<3'd1 )+$signed( -{ 2'b0,x580 }<<<3'd1 )+$signed( { 2'b0,x69 } <<<3'd1 )+$signed( -{ 3'b0,x325 }<<<3'd2)+$signed( { 1'b0,x581 }  )+$signed( -{ 1'b0,x84 } )+$signed( { 1'b0,x596 }  )+$signed( -{ 2'b0,x85 }<<<3'd1 )+$signed( -{ 1'b0,x341 } )+$signed( { 2'b0,x597 } <<<3'd1 )+$signed(11'd24);
assign y82=temp_y[82][11] ==1'b1 ? 5'd0 :  
        temp_y[82][8] ==1'b1 ? 5'd31 : 
        temp_y[82][2]==1'b1 ? temp_y[82][7:3]+1'b1 : temp_y[82][7:3];
assign temp_y[146] = 
+$signed( { 2'b0,x68 } <<<3'd1 )+$signed( { 2'b0,x324 } <<<3'd1 )+$signed( { 1'b0,x580 }  )+$signed( { 2'b0,x69 } <<<3'd1 )+$signed( -{ 1'b0,x325 } )+$signed( { 1'b0,x581 }  )+$signed( -{ 2'b0,x84 }<<<3'd1 )+$signed( -{ 2'b0,x340 }<<<3'd1 )+$signed( -{ 1'b0,x596 } )+$signed( -{ 1'b0,x85 } )+$signed( -{ 1'b0,x341 } )+$signed( -{ 1'b0,x597 } )+$signed(11'd16);
assign y146=temp_y[146][11] ==1'b1 ? 5'd0 :  
        temp_y[146][8] ==1'b1 ? 5'd31 : 
        temp_y[146][2]==1'b1 ? temp_y[146][7:3]+1'b1 : temp_y[146][7:3];
assign temp_y[210] = 
+$signed( { 1'b0,x68 }  )+$signed( -{ 1'b0,x324 } )+$signed( { 1'b0,x69 }  )+$signed( -{ 1'b0,x325 } )+$signed( { 2'b0,x84 } <<<3'd1 )+$signed( -{ 1'b0,x340 } )+$signed( -{ 1'b0,x596 } )+$signed( { 2'b0,x85 } <<<3'd1 )+$signed( -{ 1'b0,x341 } )+$signed( -{ 2'b0,x597 }<<<3'd1 )+$signed(11'd40);
assign y210=temp_y[210][11] ==1'b1 ? 5'd0 :  
        temp_y[210][8] ==1'b1 ? 5'd31 : 
        temp_y[210][2]==1'b1 ? temp_y[210][7:3]+1'b1 : temp_y[210][7:3];
assign temp_y[274] = 
+$signed( -{ 1'b0,x68 } )+$signed( { 2'b0,x324 } <<<3'd1 )+$signed( -{ 1'b0,x580 } )+$signed( -{ 1'b0,x69 } )+$signed( { 2'b0,x325 } <<<3'd1 )+$signed( -{ 2'b0,x581 }<<<3'd1 )+$signed( -{ 1'b0,x84 } )+$signed( { 2'b0,x340 } <<<3'd1 )+$signed( -{ 1'b0,x596 } )+$signed( -{ 2'b0,x85 }<<<3'd1 )+$signed( { 3'b0,x341 }<<<3'd2 )+$signed( -{ 2'b0,x597 }<<<3'd1 )+$signed(11'd32);
assign y274=temp_y[274][11] ==1'b1 ? 5'd0 :  
        temp_y[274][8] ==1'b1 ? 5'd31 : 
        temp_y[274][2]==1'b1 ? temp_y[274][7:3]+1'b1 : temp_y[274][7:3];
assign temp_y[338] = 
+$signed( -{ 1'b0,x68 } )+$signed( -{ 2'b0,x324 }<<<3'd1 )+$signed( -{ 1'b0,x580 } )+$signed( { 1'b0,x69 }  )+$signed( { 2'b0,x325 } <<<3'd1 )+$signed( { 1'b0,x581 }  )+$signed( { 1'b0,x84 }  )+$signed( { 2'b0,x340 } <<<3'd1 )+$signed( { 2'b0,x596 } <<<3'd1 )+$signed( -{ 1'b0,x85 } )+$signed( -{ 2'b0,x341 }<<<3'd1 )+$signed( -{ 1'b0,x597 } )-$signed(11'd68);
assign y338=temp_y[338][11] ==1'b1 ? 5'd0 :  
        temp_y[338][8] ==1'b1 ? 5'd31 : 
        temp_y[338][2]==1'b1 ? temp_y[338][7:3]+1'b1 : temp_y[338][7:3];
assign temp_y[402] = 
+$signed( { 1'b0,x324 }  )+$signed( { 1'b0,x581 }  )+$signed( { 1'b0,x597 }  )-$signed(11'd108);
assign y402=temp_y[402][11] ==1'b1 ? 5'd0 :  
        temp_y[402][8] ==1'b1 ? 5'd31 : 
        temp_y[402][2]==1'b1 ? temp_y[402][7:3]+1'b1 : temp_y[402][7:3];
assign temp_y[466] = 
+$signed( -{ 2'b0,x68 }<<<3'd1 )+$signed( { 2'b0,x580 } <<<3'd1 )+$signed( -{ 2'b0,x69 }<<<3'd1 )+$signed( { 1'b0,x325 }  )+$signed( { 1'b0,x581 }  )+$signed( -{ 2'b0,x84 }<<<3'd1 )+$signed( { 1'b0,x340 }  )+$signed( { 1'b0,x596 }  )+$signed( -{ 1'b0,x85 } )+$signed(11'd64);
assign y466=temp_y[466][11] ==1'b1 ? 5'd0 :  
        temp_y[466][8] ==1'b1 ? 5'd31 : 
        temp_y[466][2]==1'b1 ? temp_y[466][7:3]+1'b1 : temp_y[466][7:3];
assign temp_y[530] = 
+$signed( -{ 2'b0,x68 }<<<3'd1 )+$signed( -{ 1'b0,x324 } )+$signed( -{ 3'b0,x69 }<<<3'd2)+$signed( { 1'b0,x84 }  )+$signed( { 1'b0,x340 }  )+$signed( { 3'b0,x85 }<<<3'd2 )+$signed(11'd16);
assign y530=temp_y[530][11] ==1'b1 ? 5'd0 :  
        temp_y[530][8] ==1'b1 ? 5'd31 : 
        temp_y[530][2]==1'b1 ? temp_y[530][7:3]+1'b1 : temp_y[530][7:3];
assign temp_y[594] = 
+$signed( { 2'b0,x324 } <<<3'd1 )+$signed( { 2'b0,x580 } <<<3'd1 )+$signed( -{ 1'b0,x69 } )+$signed( -{ 2'b0,x325 }<<<3'd1 )+$signed( -{ 2'b0,x581 }<<<3'd1 )+$signed( { 2'b0,x340 } <<<3'd1 )+$signed( { 1'b0,x596 }  )+$signed( -{ 2'b0,x341 }<<<3'd1 )-$signed(11'd8);
assign y594=temp_y[594][11] ==1'b1 ? 5'd0 :  
        temp_y[594][8] ==1'b1 ? 5'd31 : 
        temp_y[594][2]==1'b1 ? temp_y[594][7:3]+1'b1 : temp_y[594][7:3];
assign temp_y[19] = 
+$signed( -{ 2'b0,x326 }<<<3'd1 )+$signed( -{ 1'b0,x582 } )+$signed( { 1'b0,x71 }  )+$signed( { 1'b0,x327 }  )+$signed( { 1'b0,x583 }  )+$signed( -{ 2'b0,x342 }<<<3'd1 )+$signed( -{ 2'b0,x598 }<<<3'd1 )+$signed( { 2'b0,x343 } <<<3'd1 )+$signed( { 2'b0,x599 } <<<3'd1 )-$signed(11'd16);
assign y19=temp_y[19][11] ==1'b1 ? 5'd0 :  
        temp_y[19][8] ==1'b1 ? 5'd31 : 
        temp_y[19][2]==1'b1 ? temp_y[19][7:3]+1'b1 : temp_y[19][7:3];
assign temp_y[83] = 
+$signed( { 3'b0,x70 }<<<3'd2 )+$signed( -{ 2'b0,x326 }<<<3'd1 )+$signed( -{ 2'b0,x582 }<<<3'd1 )+$signed( { 2'b0,x71 } <<<3'd1 )+$signed( -{ 3'b0,x327 }<<<3'd2)+$signed( { 1'b0,x583 }  )+$signed( -{ 1'b0,x86 } )+$signed( { 1'b0,x598 }  )+$signed( -{ 2'b0,x87 }<<<3'd1 )+$signed( -{ 1'b0,x343 } )+$signed( { 2'b0,x599 } <<<3'd1 )+$signed(11'd24);
assign y83=temp_y[83][11] ==1'b1 ? 5'd0 :  
        temp_y[83][8] ==1'b1 ? 5'd31 : 
        temp_y[83][2]==1'b1 ? temp_y[83][7:3]+1'b1 : temp_y[83][7:3];
assign temp_y[147] = 
+$signed( { 2'b0,x70 } <<<3'd1 )+$signed( { 2'b0,x326 } <<<3'd1 )+$signed( { 1'b0,x582 }  )+$signed( { 2'b0,x71 } <<<3'd1 )+$signed( -{ 1'b0,x327 } )+$signed( { 1'b0,x583 }  )+$signed( -{ 2'b0,x86 }<<<3'd1 )+$signed( -{ 2'b0,x342 }<<<3'd1 )+$signed( -{ 1'b0,x598 } )+$signed( -{ 1'b0,x87 } )+$signed( -{ 1'b0,x343 } )+$signed( -{ 1'b0,x599 } )+$signed(11'd16);
assign y147=temp_y[147][11] ==1'b1 ? 5'd0 :  
        temp_y[147][8] ==1'b1 ? 5'd31 : 
        temp_y[147][2]==1'b1 ? temp_y[147][7:3]+1'b1 : temp_y[147][7:3];
assign temp_y[211] = 
+$signed( { 1'b0,x70 }  )+$signed( -{ 1'b0,x326 } )+$signed( { 1'b0,x71 }  )+$signed( -{ 1'b0,x327 } )+$signed( { 2'b0,x86 } <<<3'd1 )+$signed( -{ 1'b0,x342 } )+$signed( -{ 1'b0,x598 } )+$signed( { 2'b0,x87 } <<<3'd1 )+$signed( -{ 1'b0,x343 } )+$signed( -{ 2'b0,x599 }<<<3'd1 )+$signed(11'd40);
assign y211=temp_y[211][11] ==1'b1 ? 5'd0 :  
        temp_y[211][8] ==1'b1 ? 5'd31 : 
        temp_y[211][2]==1'b1 ? temp_y[211][7:3]+1'b1 : temp_y[211][7:3];
assign temp_y[275] = 
+$signed( -{ 1'b0,x70 } )+$signed( { 2'b0,x326 } <<<3'd1 )+$signed( -{ 1'b0,x582 } )+$signed( -{ 1'b0,x71 } )+$signed( { 2'b0,x327 } <<<3'd1 )+$signed( -{ 2'b0,x583 }<<<3'd1 )+$signed( -{ 1'b0,x86 } )+$signed( { 2'b0,x342 } <<<3'd1 )+$signed( -{ 1'b0,x598 } )+$signed( -{ 2'b0,x87 }<<<3'd1 )+$signed( { 3'b0,x343 }<<<3'd2 )+$signed( -{ 2'b0,x599 }<<<3'd1 )+$signed(11'd32);
assign y275=temp_y[275][11] ==1'b1 ? 5'd0 :  
        temp_y[275][8] ==1'b1 ? 5'd31 : 
        temp_y[275][2]==1'b1 ? temp_y[275][7:3]+1'b1 : temp_y[275][7:3];
assign temp_y[339] = 
+$signed( -{ 1'b0,x70 } )+$signed( -{ 2'b0,x326 }<<<3'd1 )+$signed( -{ 1'b0,x582 } )+$signed( { 1'b0,x71 }  )+$signed( { 2'b0,x327 } <<<3'd1 )+$signed( { 1'b0,x583 }  )+$signed( { 1'b0,x86 }  )+$signed( { 2'b0,x342 } <<<3'd1 )+$signed( { 2'b0,x598 } <<<3'd1 )+$signed( -{ 1'b0,x87 } )+$signed( -{ 2'b0,x343 }<<<3'd1 )+$signed( -{ 1'b0,x599 } )-$signed(11'd68);
assign y339=temp_y[339][11] ==1'b1 ? 5'd0 :  
        temp_y[339][8] ==1'b1 ? 5'd31 : 
        temp_y[339][2]==1'b1 ? temp_y[339][7:3]+1'b1 : temp_y[339][7:3];
assign temp_y[403] = 
+$signed( { 1'b0,x326 }  )+$signed( { 1'b0,x583 }  )+$signed( { 1'b0,x599 }  )-$signed(11'd108);
assign y403=temp_y[403][11] ==1'b1 ? 5'd0 :  
        temp_y[403][8] ==1'b1 ? 5'd31 : 
        temp_y[403][2]==1'b1 ? temp_y[403][7:3]+1'b1 : temp_y[403][7:3];
assign temp_y[467] = 
+$signed( -{ 2'b0,x70 }<<<3'd1 )+$signed( { 2'b0,x582 } <<<3'd1 )+$signed( -{ 2'b0,x71 }<<<3'd1 )+$signed( { 1'b0,x327 }  )+$signed( { 1'b0,x583 }  )+$signed( -{ 2'b0,x86 }<<<3'd1 )+$signed( { 1'b0,x342 }  )+$signed( { 1'b0,x598 }  )+$signed( -{ 1'b0,x87 } )+$signed(11'd64);
assign y467=temp_y[467][11] ==1'b1 ? 5'd0 :  
        temp_y[467][8] ==1'b1 ? 5'd31 : 
        temp_y[467][2]==1'b1 ? temp_y[467][7:3]+1'b1 : temp_y[467][7:3];
assign temp_y[531] = 
+$signed( -{ 2'b0,x70 }<<<3'd1 )+$signed( -{ 1'b0,x326 } )+$signed( -{ 3'b0,x71 }<<<3'd2)+$signed( { 1'b0,x86 }  )+$signed( { 1'b0,x342 }  )+$signed( { 3'b0,x87 }<<<3'd2 )+$signed(11'd16);
assign y531=temp_y[531][11] ==1'b1 ? 5'd0 :  
        temp_y[531][8] ==1'b1 ? 5'd31 : 
        temp_y[531][2]==1'b1 ? temp_y[531][7:3]+1'b1 : temp_y[531][7:3];
assign temp_y[595] = 
+$signed( { 2'b0,x326 } <<<3'd1 )+$signed( { 2'b0,x582 } <<<3'd1 )+$signed( -{ 1'b0,x71 } )+$signed( -{ 2'b0,x327 }<<<3'd1 )+$signed( -{ 2'b0,x583 }<<<3'd1 )+$signed( { 2'b0,x342 } <<<3'd1 )+$signed( { 1'b0,x598 }  )+$signed( -{ 2'b0,x343 }<<<3'd1 )-$signed(11'd8);
assign y595=temp_y[595][11] ==1'b1 ? 5'd0 :  
        temp_y[595][8] ==1'b1 ? 5'd31 : 
        temp_y[595][2]==1'b1 ? temp_y[595][7:3]+1'b1 : temp_y[595][7:3];
assign temp_y[20] = 
+$signed( -{ 2'b0,x328 }<<<3'd1 )+$signed( -{ 1'b0,x584 } )+$signed( { 1'b0,x73 }  )+$signed( { 1'b0,x329 }  )+$signed( { 1'b0,x585 }  )+$signed( -{ 2'b0,x344 }<<<3'd1 )+$signed( -{ 2'b0,x600 }<<<3'd1 )+$signed( { 2'b0,x345 } <<<3'd1 )+$signed( { 2'b0,x601 } <<<3'd1 )-$signed(11'd16);
assign y20=temp_y[20][11] ==1'b1 ? 5'd0 :  
        temp_y[20][8] ==1'b1 ? 5'd31 : 
        temp_y[20][2]==1'b1 ? temp_y[20][7:3]+1'b1 : temp_y[20][7:3];
assign temp_y[84] = 
+$signed( { 3'b0,x72 }<<<3'd2 )+$signed( -{ 2'b0,x328 }<<<3'd1 )+$signed( -{ 2'b0,x584 }<<<3'd1 )+$signed( { 2'b0,x73 } <<<3'd1 )+$signed( -{ 3'b0,x329 }<<<3'd2)+$signed( { 1'b0,x585 }  )+$signed( -{ 1'b0,x88 } )+$signed( { 1'b0,x600 }  )+$signed( -{ 2'b0,x89 }<<<3'd1 )+$signed( -{ 1'b0,x345 } )+$signed( { 2'b0,x601 } <<<3'd1 )+$signed(11'd24);
assign y84=temp_y[84][11] ==1'b1 ? 5'd0 :  
        temp_y[84][8] ==1'b1 ? 5'd31 : 
        temp_y[84][2]==1'b1 ? temp_y[84][7:3]+1'b1 : temp_y[84][7:3];
assign temp_y[148] = 
+$signed( { 2'b0,x72 } <<<3'd1 )+$signed( { 2'b0,x328 } <<<3'd1 )+$signed( { 1'b0,x584 }  )+$signed( { 2'b0,x73 } <<<3'd1 )+$signed( -{ 1'b0,x329 } )+$signed( { 1'b0,x585 }  )+$signed( -{ 2'b0,x88 }<<<3'd1 )+$signed( -{ 2'b0,x344 }<<<3'd1 )+$signed( -{ 1'b0,x600 } )+$signed( -{ 1'b0,x89 } )+$signed( -{ 1'b0,x345 } )+$signed( -{ 1'b0,x601 } )+$signed(11'd16);
assign y148=temp_y[148][11] ==1'b1 ? 5'd0 :  
        temp_y[148][8] ==1'b1 ? 5'd31 : 
        temp_y[148][2]==1'b1 ? temp_y[148][7:3]+1'b1 : temp_y[148][7:3];
assign temp_y[212] = 
+$signed( { 1'b0,x72 }  )+$signed( -{ 1'b0,x328 } )+$signed( { 1'b0,x73 }  )+$signed( -{ 1'b0,x329 } )+$signed( { 2'b0,x88 } <<<3'd1 )+$signed( -{ 1'b0,x344 } )+$signed( -{ 1'b0,x600 } )+$signed( { 2'b0,x89 } <<<3'd1 )+$signed( -{ 1'b0,x345 } )+$signed( -{ 2'b0,x601 }<<<3'd1 )+$signed(11'd40);
assign y212=temp_y[212][11] ==1'b1 ? 5'd0 :  
        temp_y[212][8] ==1'b1 ? 5'd31 : 
        temp_y[212][2]==1'b1 ? temp_y[212][7:3]+1'b1 : temp_y[212][7:3];
assign temp_y[276] = 
+$signed( -{ 1'b0,x72 } )+$signed( { 2'b0,x328 } <<<3'd1 )+$signed( -{ 1'b0,x584 } )+$signed( -{ 1'b0,x73 } )+$signed( { 2'b0,x329 } <<<3'd1 )+$signed( -{ 2'b0,x585 }<<<3'd1 )+$signed( -{ 1'b0,x88 } )+$signed( { 2'b0,x344 } <<<3'd1 )+$signed( -{ 1'b0,x600 } )+$signed( -{ 2'b0,x89 }<<<3'd1 )+$signed( { 3'b0,x345 }<<<3'd2 )+$signed( -{ 2'b0,x601 }<<<3'd1 )+$signed(11'd32);
assign y276=temp_y[276][11] ==1'b1 ? 5'd0 :  
        temp_y[276][8] ==1'b1 ? 5'd31 : 
        temp_y[276][2]==1'b1 ? temp_y[276][7:3]+1'b1 : temp_y[276][7:3];
assign temp_y[340] = 
+$signed( -{ 1'b0,x72 } )+$signed( -{ 2'b0,x328 }<<<3'd1 )+$signed( -{ 1'b0,x584 } )+$signed( { 1'b0,x73 }  )+$signed( { 2'b0,x329 } <<<3'd1 )+$signed( { 1'b0,x585 }  )+$signed( { 1'b0,x88 }  )+$signed( { 2'b0,x344 } <<<3'd1 )+$signed( { 2'b0,x600 } <<<3'd1 )+$signed( -{ 1'b0,x89 } )+$signed( -{ 2'b0,x345 }<<<3'd1 )+$signed( -{ 1'b0,x601 } )-$signed(11'd68);
assign y340=temp_y[340][11] ==1'b1 ? 5'd0 :  
        temp_y[340][8] ==1'b1 ? 5'd31 : 
        temp_y[340][2]==1'b1 ? temp_y[340][7:3]+1'b1 : temp_y[340][7:3];
assign temp_y[404] = 
+$signed( { 1'b0,x328 }  )+$signed( { 1'b0,x585 }  )+$signed( { 1'b0,x601 }  )-$signed(11'd108);
assign y404=temp_y[404][11] ==1'b1 ? 5'd0 :  
        temp_y[404][8] ==1'b1 ? 5'd31 : 
        temp_y[404][2]==1'b1 ? temp_y[404][7:3]+1'b1 : temp_y[404][7:3];
assign temp_y[468] = 
+$signed( -{ 2'b0,x72 }<<<3'd1 )+$signed( { 2'b0,x584 } <<<3'd1 )+$signed( -{ 2'b0,x73 }<<<3'd1 )+$signed( { 1'b0,x329 }  )+$signed( { 1'b0,x585 }  )+$signed( -{ 2'b0,x88 }<<<3'd1 )+$signed( { 1'b0,x344 }  )+$signed( { 1'b0,x600 }  )+$signed( -{ 1'b0,x89 } )+$signed(11'd64);
assign y468=temp_y[468][11] ==1'b1 ? 5'd0 :  
        temp_y[468][8] ==1'b1 ? 5'd31 : 
        temp_y[468][2]==1'b1 ? temp_y[468][7:3]+1'b1 : temp_y[468][7:3];
assign temp_y[532] = 
+$signed( -{ 2'b0,x72 }<<<3'd1 )+$signed( -{ 1'b0,x328 } )+$signed( -{ 3'b0,x73 }<<<3'd2)+$signed( { 1'b0,x88 }  )+$signed( { 1'b0,x344 }  )+$signed( { 3'b0,x89 }<<<3'd2 )+$signed(11'd16);
assign y532=temp_y[532][11] ==1'b1 ? 5'd0 :  
        temp_y[532][8] ==1'b1 ? 5'd31 : 
        temp_y[532][2]==1'b1 ? temp_y[532][7:3]+1'b1 : temp_y[532][7:3];
assign temp_y[596] = 
+$signed( { 2'b0,x328 } <<<3'd1 )+$signed( { 2'b0,x584 } <<<3'd1 )+$signed( -{ 1'b0,x73 } )+$signed( -{ 2'b0,x329 }<<<3'd1 )+$signed( -{ 2'b0,x585 }<<<3'd1 )+$signed( { 2'b0,x344 } <<<3'd1 )+$signed( { 1'b0,x600 }  )+$signed( -{ 2'b0,x345 }<<<3'd1 )-$signed(11'd8);
assign y596=temp_y[596][11] ==1'b1 ? 5'd0 :  
        temp_y[596][8] ==1'b1 ? 5'd31 : 
        temp_y[596][2]==1'b1 ? temp_y[596][7:3]+1'b1 : temp_y[596][7:3];
assign temp_y[21] = 
+$signed( -{ 2'b0,x330 }<<<3'd1 )+$signed( -{ 1'b0,x586 } )+$signed( { 1'b0,x75 }  )+$signed( { 1'b0,x331 }  )+$signed( { 1'b0,x587 }  )+$signed( -{ 2'b0,x346 }<<<3'd1 )+$signed( -{ 2'b0,x602 }<<<3'd1 )+$signed( { 2'b0,x347 } <<<3'd1 )+$signed( { 2'b0,x603 } <<<3'd1 )-$signed(11'd16);
assign y21=temp_y[21][11] ==1'b1 ? 5'd0 :  
        temp_y[21][8] ==1'b1 ? 5'd31 : 
        temp_y[21][2]==1'b1 ? temp_y[21][7:3]+1'b1 : temp_y[21][7:3];
assign temp_y[85] = 
+$signed( { 3'b0,x74 }<<<3'd2 )+$signed( -{ 2'b0,x330 }<<<3'd1 )+$signed( -{ 2'b0,x586 }<<<3'd1 )+$signed( { 2'b0,x75 } <<<3'd1 )+$signed( -{ 3'b0,x331 }<<<3'd2)+$signed( { 1'b0,x587 }  )+$signed( -{ 1'b0,x90 } )+$signed( { 1'b0,x602 }  )+$signed( -{ 2'b0,x91 }<<<3'd1 )+$signed( -{ 1'b0,x347 } )+$signed( { 2'b0,x603 } <<<3'd1 )+$signed(11'd24);
assign y85=temp_y[85][11] ==1'b1 ? 5'd0 :  
        temp_y[85][8] ==1'b1 ? 5'd31 : 
        temp_y[85][2]==1'b1 ? temp_y[85][7:3]+1'b1 : temp_y[85][7:3];
assign temp_y[149] = 
+$signed( { 2'b0,x74 } <<<3'd1 )+$signed( { 2'b0,x330 } <<<3'd1 )+$signed( { 1'b0,x586 }  )+$signed( { 2'b0,x75 } <<<3'd1 )+$signed( -{ 1'b0,x331 } )+$signed( { 1'b0,x587 }  )+$signed( -{ 2'b0,x90 }<<<3'd1 )+$signed( -{ 2'b0,x346 }<<<3'd1 )+$signed( -{ 1'b0,x602 } )+$signed( -{ 1'b0,x91 } )+$signed( -{ 1'b0,x347 } )+$signed( -{ 1'b0,x603 } )+$signed(11'd16);
assign y149=temp_y[149][11] ==1'b1 ? 5'd0 :  
        temp_y[149][8] ==1'b1 ? 5'd31 : 
        temp_y[149][2]==1'b1 ? temp_y[149][7:3]+1'b1 : temp_y[149][7:3];
assign temp_y[213] = 
+$signed( { 1'b0,x74 }  )+$signed( -{ 1'b0,x330 } )+$signed( { 1'b0,x75 }  )+$signed( -{ 1'b0,x331 } )+$signed( { 2'b0,x90 } <<<3'd1 )+$signed( -{ 1'b0,x346 } )+$signed( -{ 1'b0,x602 } )+$signed( { 2'b0,x91 } <<<3'd1 )+$signed( -{ 1'b0,x347 } )+$signed( -{ 2'b0,x603 }<<<3'd1 )+$signed(11'd40);
assign y213=temp_y[213][11] ==1'b1 ? 5'd0 :  
        temp_y[213][8] ==1'b1 ? 5'd31 : 
        temp_y[213][2]==1'b1 ? temp_y[213][7:3]+1'b1 : temp_y[213][7:3];
assign temp_y[277] = 
+$signed( -{ 1'b0,x74 } )+$signed( { 2'b0,x330 } <<<3'd1 )+$signed( -{ 1'b0,x586 } )+$signed( -{ 1'b0,x75 } )+$signed( { 2'b0,x331 } <<<3'd1 )+$signed( -{ 2'b0,x587 }<<<3'd1 )+$signed( -{ 1'b0,x90 } )+$signed( { 2'b0,x346 } <<<3'd1 )+$signed( -{ 1'b0,x602 } )+$signed( -{ 2'b0,x91 }<<<3'd1 )+$signed( { 3'b0,x347 }<<<3'd2 )+$signed( -{ 2'b0,x603 }<<<3'd1 )+$signed(11'd32);
assign y277=temp_y[277][11] ==1'b1 ? 5'd0 :  
        temp_y[277][8] ==1'b1 ? 5'd31 : 
        temp_y[277][2]==1'b1 ? temp_y[277][7:3]+1'b1 : temp_y[277][7:3];
assign temp_y[341] = 
+$signed( -{ 1'b0,x74 } )+$signed( -{ 2'b0,x330 }<<<3'd1 )+$signed( -{ 1'b0,x586 } )+$signed( { 1'b0,x75 }  )+$signed( { 2'b0,x331 } <<<3'd1 )+$signed( { 1'b0,x587 }  )+$signed( { 1'b0,x90 }  )+$signed( { 2'b0,x346 } <<<3'd1 )+$signed( { 2'b0,x602 } <<<3'd1 )+$signed( -{ 1'b0,x91 } )+$signed( -{ 2'b0,x347 }<<<3'd1 )+$signed( -{ 1'b0,x603 } )-$signed(11'd68);
assign y341=temp_y[341][11] ==1'b1 ? 5'd0 :  
        temp_y[341][8] ==1'b1 ? 5'd31 : 
        temp_y[341][2]==1'b1 ? temp_y[341][7:3]+1'b1 : temp_y[341][7:3];
assign temp_y[405] = 
+$signed( { 1'b0,x330 }  )+$signed( { 1'b0,x587 }  )+$signed( { 1'b0,x603 }  )-$signed(11'd108);
assign y405=temp_y[405][11] ==1'b1 ? 5'd0 :  
        temp_y[405][8] ==1'b1 ? 5'd31 : 
        temp_y[405][2]==1'b1 ? temp_y[405][7:3]+1'b1 : temp_y[405][7:3];
assign temp_y[469] = 
+$signed( -{ 2'b0,x74 }<<<3'd1 )+$signed( { 2'b0,x586 } <<<3'd1 )+$signed( -{ 2'b0,x75 }<<<3'd1 )+$signed( { 1'b0,x331 }  )+$signed( { 1'b0,x587 }  )+$signed( -{ 2'b0,x90 }<<<3'd1 )+$signed( { 1'b0,x346 }  )+$signed( { 1'b0,x602 }  )+$signed( -{ 1'b0,x91 } )+$signed(11'd64);
assign y469=temp_y[469][11] ==1'b1 ? 5'd0 :  
        temp_y[469][8] ==1'b1 ? 5'd31 : 
        temp_y[469][2]==1'b1 ? temp_y[469][7:3]+1'b1 : temp_y[469][7:3];
assign temp_y[533] = 
+$signed( -{ 2'b0,x74 }<<<3'd1 )+$signed( -{ 1'b0,x330 } )+$signed( -{ 3'b0,x75 }<<<3'd2)+$signed( { 1'b0,x90 }  )+$signed( { 1'b0,x346 }  )+$signed( { 3'b0,x91 }<<<3'd2 )+$signed(11'd16);
assign y533=temp_y[533][11] ==1'b1 ? 5'd0 :  
        temp_y[533][8] ==1'b1 ? 5'd31 : 
        temp_y[533][2]==1'b1 ? temp_y[533][7:3]+1'b1 : temp_y[533][7:3];
assign temp_y[597] = 
+$signed( { 2'b0,x330 } <<<3'd1 )+$signed( { 2'b0,x586 } <<<3'd1 )+$signed( -{ 1'b0,x75 } )+$signed( -{ 2'b0,x331 }<<<3'd1 )+$signed( -{ 2'b0,x587 }<<<3'd1 )+$signed( { 2'b0,x346 } <<<3'd1 )+$signed( { 1'b0,x602 }  )+$signed( -{ 2'b0,x347 }<<<3'd1 )-$signed(11'd8);
assign y597=temp_y[597][11] ==1'b1 ? 5'd0 :  
        temp_y[597][8] ==1'b1 ? 5'd31 : 
        temp_y[597][2]==1'b1 ? temp_y[597][7:3]+1'b1 : temp_y[597][7:3];
assign temp_y[22] = 
+$signed( -{ 2'b0,x332 }<<<3'd1 )+$signed( -{ 1'b0,x588 } )+$signed( { 1'b0,x77 }  )+$signed( { 1'b0,x333 }  )+$signed( { 1'b0,x589 }  )+$signed( -{ 2'b0,x348 }<<<3'd1 )+$signed( -{ 2'b0,x604 }<<<3'd1 )+$signed( { 2'b0,x349 } <<<3'd1 )+$signed( { 2'b0,x605 } <<<3'd1 )-$signed(11'd16);
assign y22=temp_y[22][11] ==1'b1 ? 5'd0 :  
        temp_y[22][8] ==1'b1 ? 5'd31 : 
        temp_y[22][2]==1'b1 ? temp_y[22][7:3]+1'b1 : temp_y[22][7:3];
assign temp_y[86] = 
+$signed( { 3'b0,x76 }<<<3'd2 )+$signed( -{ 2'b0,x332 }<<<3'd1 )+$signed( -{ 2'b0,x588 }<<<3'd1 )+$signed( { 2'b0,x77 } <<<3'd1 )+$signed( -{ 3'b0,x333 }<<<3'd2)+$signed( { 1'b0,x589 }  )+$signed( -{ 1'b0,x92 } )+$signed( { 1'b0,x604 }  )+$signed( -{ 2'b0,x93 }<<<3'd1 )+$signed( -{ 1'b0,x349 } )+$signed( { 2'b0,x605 } <<<3'd1 )+$signed(11'd24);
assign y86=temp_y[86][11] ==1'b1 ? 5'd0 :  
        temp_y[86][8] ==1'b1 ? 5'd31 : 
        temp_y[86][2]==1'b1 ? temp_y[86][7:3]+1'b1 : temp_y[86][7:3];
assign temp_y[150] = 
+$signed( { 2'b0,x76 } <<<3'd1 )+$signed( { 2'b0,x332 } <<<3'd1 )+$signed( { 1'b0,x588 }  )+$signed( { 2'b0,x77 } <<<3'd1 )+$signed( -{ 1'b0,x333 } )+$signed( { 1'b0,x589 }  )+$signed( -{ 2'b0,x92 }<<<3'd1 )+$signed( -{ 2'b0,x348 }<<<3'd1 )+$signed( -{ 1'b0,x604 } )+$signed( -{ 1'b0,x93 } )+$signed( -{ 1'b0,x349 } )+$signed( -{ 1'b0,x605 } )+$signed(11'd16);
assign y150=temp_y[150][11] ==1'b1 ? 5'd0 :  
        temp_y[150][8] ==1'b1 ? 5'd31 : 
        temp_y[150][2]==1'b1 ? temp_y[150][7:3]+1'b1 : temp_y[150][7:3];
assign temp_y[214] = 
+$signed( { 1'b0,x76 }  )+$signed( -{ 1'b0,x332 } )+$signed( { 1'b0,x77 }  )+$signed( -{ 1'b0,x333 } )+$signed( { 2'b0,x92 } <<<3'd1 )+$signed( -{ 1'b0,x348 } )+$signed( -{ 1'b0,x604 } )+$signed( { 2'b0,x93 } <<<3'd1 )+$signed( -{ 1'b0,x349 } )+$signed( -{ 2'b0,x605 }<<<3'd1 )+$signed(11'd40);
assign y214=temp_y[214][11] ==1'b1 ? 5'd0 :  
        temp_y[214][8] ==1'b1 ? 5'd31 : 
        temp_y[214][2]==1'b1 ? temp_y[214][7:3]+1'b1 : temp_y[214][7:3];
assign temp_y[278] = 
+$signed( -{ 1'b0,x76 } )+$signed( { 2'b0,x332 } <<<3'd1 )+$signed( -{ 1'b0,x588 } )+$signed( -{ 1'b0,x77 } )+$signed( { 2'b0,x333 } <<<3'd1 )+$signed( -{ 2'b0,x589 }<<<3'd1 )+$signed( -{ 1'b0,x92 } )+$signed( { 2'b0,x348 } <<<3'd1 )+$signed( -{ 1'b0,x604 } )+$signed( -{ 2'b0,x93 }<<<3'd1 )+$signed( { 3'b0,x349 }<<<3'd2 )+$signed( -{ 2'b0,x605 }<<<3'd1 )+$signed(11'd32);
assign y278=temp_y[278][11] ==1'b1 ? 5'd0 :  
        temp_y[278][8] ==1'b1 ? 5'd31 : 
        temp_y[278][2]==1'b1 ? temp_y[278][7:3]+1'b1 : temp_y[278][7:3];
assign temp_y[342] = 
+$signed( -{ 1'b0,x76 } )+$signed( -{ 2'b0,x332 }<<<3'd1 )+$signed( -{ 1'b0,x588 } )+$signed( { 1'b0,x77 }  )+$signed( { 2'b0,x333 } <<<3'd1 )+$signed( { 1'b0,x589 }  )+$signed( { 1'b0,x92 }  )+$signed( { 2'b0,x348 } <<<3'd1 )+$signed( { 2'b0,x604 } <<<3'd1 )+$signed( -{ 1'b0,x93 } )+$signed( -{ 2'b0,x349 }<<<3'd1 )+$signed( -{ 1'b0,x605 } )-$signed(11'd68);
assign y342=temp_y[342][11] ==1'b1 ? 5'd0 :  
        temp_y[342][8] ==1'b1 ? 5'd31 : 
        temp_y[342][2]==1'b1 ? temp_y[342][7:3]+1'b1 : temp_y[342][7:3];
assign temp_y[406] = 
+$signed( { 1'b0,x332 }  )+$signed( { 1'b0,x589 }  )+$signed( { 1'b0,x605 }  )-$signed(11'd108);
assign y406=temp_y[406][11] ==1'b1 ? 5'd0 :  
        temp_y[406][8] ==1'b1 ? 5'd31 : 
        temp_y[406][2]==1'b1 ? temp_y[406][7:3]+1'b1 : temp_y[406][7:3];
assign temp_y[470] = 
+$signed( -{ 2'b0,x76 }<<<3'd1 )+$signed( { 2'b0,x588 } <<<3'd1 )+$signed( -{ 2'b0,x77 }<<<3'd1 )+$signed( { 1'b0,x333 }  )+$signed( { 1'b0,x589 }  )+$signed( -{ 2'b0,x92 }<<<3'd1 )+$signed( { 1'b0,x348 }  )+$signed( { 1'b0,x604 }  )+$signed( -{ 1'b0,x93 } )+$signed(11'd64);
assign y470=temp_y[470][11] ==1'b1 ? 5'd0 :  
        temp_y[470][8] ==1'b1 ? 5'd31 : 
        temp_y[470][2]==1'b1 ? temp_y[470][7:3]+1'b1 : temp_y[470][7:3];
assign temp_y[534] = 
+$signed( -{ 2'b0,x76 }<<<3'd1 )+$signed( -{ 1'b0,x332 } )+$signed( -{ 3'b0,x77 }<<<3'd2)+$signed( { 1'b0,x92 }  )+$signed( { 1'b0,x348 }  )+$signed( { 3'b0,x93 }<<<3'd2 )+$signed(11'd16);
assign y534=temp_y[534][11] ==1'b1 ? 5'd0 :  
        temp_y[534][8] ==1'b1 ? 5'd31 : 
        temp_y[534][2]==1'b1 ? temp_y[534][7:3]+1'b1 : temp_y[534][7:3];
assign temp_y[598] = 
+$signed( { 2'b0,x332 } <<<3'd1 )+$signed( { 2'b0,x588 } <<<3'd1 )+$signed( -{ 1'b0,x77 } )+$signed( -{ 2'b0,x333 }<<<3'd1 )+$signed( -{ 2'b0,x589 }<<<3'd1 )+$signed( { 2'b0,x348 } <<<3'd1 )+$signed( { 1'b0,x604 }  )+$signed( -{ 2'b0,x349 }<<<3'd1 )-$signed(11'd8);
assign y598=temp_y[598][11] ==1'b1 ? 5'd0 :  
        temp_y[598][8] ==1'b1 ? 5'd31 : 
        temp_y[598][2]==1'b1 ? temp_y[598][7:3]+1'b1 : temp_y[598][7:3];
assign temp_y[23] = 
+$signed( -{ 2'b0,x334 }<<<3'd1 )+$signed( -{ 1'b0,x590 } )+$signed( { 1'b0,x79 }  )+$signed( { 1'b0,x335 }  )+$signed( { 1'b0,x591 }  )+$signed( -{ 2'b0,x350 }<<<3'd1 )+$signed( -{ 2'b0,x606 }<<<3'd1 )+$signed( { 2'b0,x351 } <<<3'd1 )+$signed( { 2'b0,x607 } <<<3'd1 )-$signed(11'd16);
assign y23=temp_y[23][11] ==1'b1 ? 5'd0 :  
        temp_y[23][8] ==1'b1 ? 5'd31 : 
        temp_y[23][2]==1'b1 ? temp_y[23][7:3]+1'b1 : temp_y[23][7:3];
assign temp_y[87] = 
+$signed( { 3'b0,x78 }<<<3'd2 )+$signed( -{ 2'b0,x334 }<<<3'd1 )+$signed( -{ 2'b0,x590 }<<<3'd1 )+$signed( { 2'b0,x79 } <<<3'd1 )+$signed( -{ 3'b0,x335 }<<<3'd2)+$signed( { 1'b0,x591 }  )+$signed( -{ 1'b0,x94 } )+$signed( { 1'b0,x606 }  )+$signed( -{ 2'b0,x95 }<<<3'd1 )+$signed( -{ 1'b0,x351 } )+$signed( { 2'b0,x607 } <<<3'd1 )+$signed(11'd24);
assign y87=temp_y[87][11] ==1'b1 ? 5'd0 :  
        temp_y[87][8] ==1'b1 ? 5'd31 : 
        temp_y[87][2]==1'b1 ? temp_y[87][7:3]+1'b1 : temp_y[87][7:3];
assign temp_y[151] = 
+$signed( { 2'b0,x78 } <<<3'd1 )+$signed( { 2'b0,x334 } <<<3'd1 )+$signed( { 1'b0,x590 }  )+$signed( { 2'b0,x79 } <<<3'd1 )+$signed( -{ 1'b0,x335 } )+$signed( { 1'b0,x591 }  )+$signed( -{ 2'b0,x94 }<<<3'd1 )+$signed( -{ 2'b0,x350 }<<<3'd1 )+$signed( -{ 1'b0,x606 } )+$signed( -{ 1'b0,x95 } )+$signed( -{ 1'b0,x351 } )+$signed( -{ 1'b0,x607 } )+$signed(11'd16);
assign y151=temp_y[151][11] ==1'b1 ? 5'd0 :  
        temp_y[151][8] ==1'b1 ? 5'd31 : 
        temp_y[151][2]==1'b1 ? temp_y[151][7:3]+1'b1 : temp_y[151][7:3];
assign temp_y[215] = 
+$signed( { 1'b0,x78 }  )+$signed( -{ 1'b0,x334 } )+$signed( { 1'b0,x79 }  )+$signed( -{ 1'b0,x335 } )+$signed( { 2'b0,x94 } <<<3'd1 )+$signed( -{ 1'b0,x350 } )+$signed( -{ 1'b0,x606 } )+$signed( { 2'b0,x95 } <<<3'd1 )+$signed( -{ 1'b0,x351 } )+$signed( -{ 2'b0,x607 }<<<3'd1 )+$signed(11'd40);
assign y215=temp_y[215][11] ==1'b1 ? 5'd0 :  
        temp_y[215][8] ==1'b1 ? 5'd31 : 
        temp_y[215][2]==1'b1 ? temp_y[215][7:3]+1'b1 : temp_y[215][7:3];
assign temp_y[279] = 
+$signed( -{ 1'b0,x78 } )+$signed( { 2'b0,x334 } <<<3'd1 )+$signed( -{ 1'b0,x590 } )+$signed( -{ 1'b0,x79 } )+$signed( { 2'b0,x335 } <<<3'd1 )+$signed( -{ 2'b0,x591 }<<<3'd1 )+$signed( -{ 1'b0,x94 } )+$signed( { 2'b0,x350 } <<<3'd1 )+$signed( -{ 1'b0,x606 } )+$signed( -{ 2'b0,x95 }<<<3'd1 )+$signed( { 3'b0,x351 }<<<3'd2 )+$signed( -{ 2'b0,x607 }<<<3'd1 )+$signed(11'd32);
assign y279=temp_y[279][11] ==1'b1 ? 5'd0 :  
        temp_y[279][8] ==1'b1 ? 5'd31 : 
        temp_y[279][2]==1'b1 ? temp_y[279][7:3]+1'b1 : temp_y[279][7:3];
assign temp_y[343] = 
+$signed( -{ 1'b0,x78 } )+$signed( -{ 2'b0,x334 }<<<3'd1 )+$signed( -{ 1'b0,x590 } )+$signed( { 1'b0,x79 }  )+$signed( { 2'b0,x335 } <<<3'd1 )+$signed( { 1'b0,x591 }  )+$signed( { 1'b0,x94 }  )+$signed( { 2'b0,x350 } <<<3'd1 )+$signed( { 2'b0,x606 } <<<3'd1 )+$signed( -{ 1'b0,x95 } )+$signed( -{ 2'b0,x351 }<<<3'd1 )+$signed( -{ 1'b0,x607 } )-$signed(11'd68);
assign y343=temp_y[343][11] ==1'b1 ? 5'd0 :  
        temp_y[343][8] ==1'b1 ? 5'd31 : 
        temp_y[343][2]==1'b1 ? temp_y[343][7:3]+1'b1 : temp_y[343][7:3];
assign temp_y[407] = 
+$signed( { 1'b0,x334 }  )+$signed( { 1'b0,x591 }  )+$signed( { 1'b0,x607 }  )-$signed(11'd108);
assign y407=temp_y[407][11] ==1'b1 ? 5'd0 :  
        temp_y[407][8] ==1'b1 ? 5'd31 : 
        temp_y[407][2]==1'b1 ? temp_y[407][7:3]+1'b1 : temp_y[407][7:3];
assign temp_y[471] = 
+$signed( -{ 2'b0,x78 }<<<3'd1 )+$signed( { 2'b0,x590 } <<<3'd1 )+$signed( -{ 2'b0,x79 }<<<3'd1 )+$signed( { 1'b0,x335 }  )+$signed( { 1'b0,x591 }  )+$signed( -{ 2'b0,x94 }<<<3'd1 )+$signed( { 1'b0,x350 }  )+$signed( { 1'b0,x606 }  )+$signed( -{ 1'b0,x95 } )+$signed(11'd64);
assign y471=temp_y[471][11] ==1'b1 ? 5'd0 :  
        temp_y[471][8] ==1'b1 ? 5'd31 : 
        temp_y[471][2]==1'b1 ? temp_y[471][7:3]+1'b1 : temp_y[471][7:3];
assign temp_y[535] = 
+$signed( -{ 2'b0,x78 }<<<3'd1 )+$signed( -{ 1'b0,x334 } )+$signed( -{ 3'b0,x79 }<<<3'd2)+$signed( { 1'b0,x94 }  )+$signed( { 1'b0,x350 }  )+$signed( { 3'b0,x95 }<<<3'd2 )+$signed(11'd16);
assign y535=temp_y[535][11] ==1'b1 ? 5'd0 :  
        temp_y[535][8] ==1'b1 ? 5'd31 : 
        temp_y[535][2]==1'b1 ? temp_y[535][7:3]+1'b1 : temp_y[535][7:3];
assign temp_y[599] = 
+$signed( { 2'b0,x334 } <<<3'd1 )+$signed( { 2'b0,x590 } <<<3'd1 )+$signed( -{ 1'b0,x79 } )+$signed( -{ 2'b0,x335 }<<<3'd1 )+$signed( -{ 2'b0,x591 }<<<3'd1 )+$signed( { 2'b0,x350 } <<<3'd1 )+$signed( { 1'b0,x606 }  )+$signed( -{ 2'b0,x351 }<<<3'd1 )-$signed(11'd8);
assign y599=temp_y[599][11] ==1'b1 ? 5'd0 :  
        temp_y[599][8] ==1'b1 ? 5'd31 : 
        temp_y[599][2]==1'b1 ? temp_y[599][7:3]+1'b1 : temp_y[599][7:3];
assign temp_y[24] = 
+$signed( -{ 2'b0,x352 }<<<3'd1 )+$signed( -{ 1'b0,x608 } )+$signed( { 1'b0,x97 }  )+$signed( { 1'b0,x353 }  )+$signed( { 1'b0,x609 }  )+$signed( -{ 2'b0,x368 }<<<3'd1 )+$signed( -{ 2'b0,x624 }<<<3'd1 )+$signed( { 2'b0,x369 } <<<3'd1 )+$signed( { 2'b0,x625 } <<<3'd1 )-$signed(11'd16);
assign y24=temp_y[24][11] ==1'b1 ? 5'd0 :  
        temp_y[24][8] ==1'b1 ? 5'd31 : 
        temp_y[24][2]==1'b1 ? temp_y[24][7:3]+1'b1 : temp_y[24][7:3];
assign temp_y[88] = 
+$signed( { 3'b0,x96 }<<<3'd2 )+$signed( -{ 2'b0,x352 }<<<3'd1 )+$signed( -{ 2'b0,x608 }<<<3'd1 )+$signed( { 2'b0,x97 } <<<3'd1 )+$signed( -{ 3'b0,x353 }<<<3'd2)+$signed( { 1'b0,x609 }  )+$signed( -{ 1'b0,x112 } )+$signed( { 1'b0,x624 }  )+$signed( -{ 2'b0,x113 }<<<3'd1 )+$signed( -{ 1'b0,x369 } )+$signed( { 2'b0,x625 } <<<3'd1 )+$signed(11'd24);
assign y88=temp_y[88][11] ==1'b1 ? 5'd0 :  
        temp_y[88][8] ==1'b1 ? 5'd31 : 
        temp_y[88][2]==1'b1 ? temp_y[88][7:3]+1'b1 : temp_y[88][7:3];
assign temp_y[152] = 
+$signed( { 2'b0,x96 } <<<3'd1 )+$signed( { 2'b0,x352 } <<<3'd1 )+$signed( { 1'b0,x608 }  )+$signed( { 2'b0,x97 } <<<3'd1 )+$signed( -{ 1'b0,x353 } )+$signed( { 1'b0,x609 }  )+$signed( -{ 2'b0,x112 }<<<3'd1 )+$signed( -{ 2'b0,x368 }<<<3'd1 )+$signed( -{ 1'b0,x624 } )+$signed( -{ 1'b0,x113 } )+$signed( -{ 1'b0,x369 } )+$signed( -{ 1'b0,x625 } )+$signed(11'd16);
assign y152=temp_y[152][11] ==1'b1 ? 5'd0 :  
        temp_y[152][8] ==1'b1 ? 5'd31 : 
        temp_y[152][2]==1'b1 ? temp_y[152][7:3]+1'b1 : temp_y[152][7:3];
assign temp_y[216] = 
+$signed( { 1'b0,x96 }  )+$signed( -{ 1'b0,x352 } )+$signed( { 1'b0,x97 }  )+$signed( -{ 1'b0,x353 } )+$signed( { 2'b0,x112 } <<<3'd1 )+$signed( -{ 1'b0,x368 } )+$signed( -{ 1'b0,x624 } )+$signed( { 2'b0,x113 } <<<3'd1 )+$signed( -{ 1'b0,x369 } )+$signed( -{ 2'b0,x625 }<<<3'd1 )+$signed(11'd40);
assign y216=temp_y[216][11] ==1'b1 ? 5'd0 :  
        temp_y[216][8] ==1'b1 ? 5'd31 : 
        temp_y[216][2]==1'b1 ? temp_y[216][7:3]+1'b1 : temp_y[216][7:3];
assign temp_y[280] = 
+$signed( -{ 1'b0,x96 } )+$signed( { 2'b0,x352 } <<<3'd1 )+$signed( -{ 1'b0,x608 } )+$signed( -{ 1'b0,x97 } )+$signed( { 2'b0,x353 } <<<3'd1 )+$signed( -{ 2'b0,x609 }<<<3'd1 )+$signed( -{ 1'b0,x112 } )+$signed( { 2'b0,x368 } <<<3'd1 )+$signed( -{ 1'b0,x624 } )+$signed( -{ 2'b0,x113 }<<<3'd1 )+$signed( { 3'b0,x369 }<<<3'd2 )+$signed( -{ 2'b0,x625 }<<<3'd1 )+$signed(11'd32);
assign y280=temp_y[280][11] ==1'b1 ? 5'd0 :  
        temp_y[280][8] ==1'b1 ? 5'd31 : 
        temp_y[280][2]==1'b1 ? temp_y[280][7:3]+1'b1 : temp_y[280][7:3];
assign temp_y[344] = 
+$signed( -{ 1'b0,x96 } )+$signed( -{ 2'b0,x352 }<<<3'd1 )+$signed( -{ 1'b0,x608 } )+$signed( { 1'b0,x97 }  )+$signed( { 2'b0,x353 } <<<3'd1 )+$signed( { 1'b0,x609 }  )+$signed( { 1'b0,x112 }  )+$signed( { 2'b0,x368 } <<<3'd1 )+$signed( { 2'b0,x624 } <<<3'd1 )+$signed( -{ 1'b0,x113 } )+$signed( -{ 2'b0,x369 }<<<3'd1 )+$signed( -{ 1'b0,x625 } )-$signed(11'd68);
assign y344=temp_y[344][11] ==1'b1 ? 5'd0 :  
        temp_y[344][8] ==1'b1 ? 5'd31 : 
        temp_y[344][2]==1'b1 ? temp_y[344][7:3]+1'b1 : temp_y[344][7:3];
assign temp_y[408] = 
+$signed( { 1'b0,x352 }  )+$signed( { 1'b0,x609 }  )+$signed( { 1'b0,x625 }  )-$signed(11'd108);
assign y408=temp_y[408][11] ==1'b1 ? 5'd0 :  
        temp_y[408][8] ==1'b1 ? 5'd31 : 
        temp_y[408][2]==1'b1 ? temp_y[408][7:3]+1'b1 : temp_y[408][7:3];
assign temp_y[472] = 
+$signed( -{ 2'b0,x96 }<<<3'd1 )+$signed( { 2'b0,x608 } <<<3'd1 )+$signed( -{ 2'b0,x97 }<<<3'd1 )+$signed( { 1'b0,x353 }  )+$signed( { 1'b0,x609 }  )+$signed( -{ 2'b0,x112 }<<<3'd1 )+$signed( { 1'b0,x368 }  )+$signed( { 1'b0,x624 }  )+$signed( -{ 1'b0,x113 } )+$signed(11'd64);
assign y472=temp_y[472][11] ==1'b1 ? 5'd0 :  
        temp_y[472][8] ==1'b1 ? 5'd31 : 
        temp_y[472][2]==1'b1 ? temp_y[472][7:3]+1'b1 : temp_y[472][7:3];
assign temp_y[536] = 
+$signed( -{ 2'b0,x96 }<<<3'd1 )+$signed( -{ 1'b0,x352 } )+$signed( -{ 3'b0,x97 }<<<3'd2)+$signed( { 1'b0,x112 }  )+$signed( { 1'b0,x368 }  )+$signed( { 3'b0,x113 }<<<3'd2 )+$signed(11'd16);
assign y536=temp_y[536][11] ==1'b1 ? 5'd0 :  
        temp_y[536][8] ==1'b1 ? 5'd31 : 
        temp_y[536][2]==1'b1 ? temp_y[536][7:3]+1'b1 : temp_y[536][7:3];
assign temp_y[600] = 
+$signed( { 2'b0,x352 } <<<3'd1 )+$signed( { 2'b0,x608 } <<<3'd1 )+$signed( -{ 1'b0,x97 } )+$signed( -{ 2'b0,x353 }<<<3'd1 )+$signed( -{ 2'b0,x609 }<<<3'd1 )+$signed( { 2'b0,x368 } <<<3'd1 )+$signed( { 1'b0,x624 }  )+$signed( -{ 2'b0,x369 }<<<3'd1 )-$signed(11'd8);
assign y600=temp_y[600][11] ==1'b1 ? 5'd0 :  
        temp_y[600][8] ==1'b1 ? 5'd31 : 
        temp_y[600][2]==1'b1 ? temp_y[600][7:3]+1'b1 : temp_y[600][7:3];
assign temp_y[25] = 
+$signed( -{ 2'b0,x354 }<<<3'd1 )+$signed( -{ 1'b0,x610 } )+$signed( { 1'b0,x99 }  )+$signed( { 1'b0,x355 }  )+$signed( { 1'b0,x611 }  )+$signed( -{ 2'b0,x370 }<<<3'd1 )+$signed( -{ 2'b0,x626 }<<<3'd1 )+$signed( { 2'b0,x371 } <<<3'd1 )+$signed( { 2'b0,x627 } <<<3'd1 )-$signed(11'd16);
assign y25=temp_y[25][11] ==1'b1 ? 5'd0 :  
        temp_y[25][8] ==1'b1 ? 5'd31 : 
        temp_y[25][2]==1'b1 ? temp_y[25][7:3]+1'b1 : temp_y[25][7:3];
assign temp_y[89] = 
+$signed( { 3'b0,x98 }<<<3'd2 )+$signed( -{ 2'b0,x354 }<<<3'd1 )+$signed( -{ 2'b0,x610 }<<<3'd1 )+$signed( { 2'b0,x99 } <<<3'd1 )+$signed( -{ 3'b0,x355 }<<<3'd2)+$signed( { 1'b0,x611 }  )+$signed( -{ 1'b0,x114 } )+$signed( { 1'b0,x626 }  )+$signed( -{ 2'b0,x115 }<<<3'd1 )+$signed( -{ 1'b0,x371 } )+$signed( { 2'b0,x627 } <<<3'd1 )+$signed(11'd24);
assign y89=temp_y[89][11] ==1'b1 ? 5'd0 :  
        temp_y[89][8] ==1'b1 ? 5'd31 : 
        temp_y[89][2]==1'b1 ? temp_y[89][7:3]+1'b1 : temp_y[89][7:3];
assign temp_y[153] = 
+$signed( { 2'b0,x98 } <<<3'd1 )+$signed( { 2'b0,x354 } <<<3'd1 )+$signed( { 1'b0,x610 }  )+$signed( { 2'b0,x99 } <<<3'd1 )+$signed( -{ 1'b0,x355 } )+$signed( { 1'b0,x611 }  )+$signed( -{ 2'b0,x114 }<<<3'd1 )+$signed( -{ 2'b0,x370 }<<<3'd1 )+$signed( -{ 1'b0,x626 } )+$signed( -{ 1'b0,x115 } )+$signed( -{ 1'b0,x371 } )+$signed( -{ 1'b0,x627 } )+$signed(11'd16);
assign y153=temp_y[153][11] ==1'b1 ? 5'd0 :  
        temp_y[153][8] ==1'b1 ? 5'd31 : 
        temp_y[153][2]==1'b1 ? temp_y[153][7:3]+1'b1 : temp_y[153][7:3];
assign temp_y[217] = 
+$signed( { 1'b0,x98 }  )+$signed( -{ 1'b0,x354 } )+$signed( { 1'b0,x99 }  )+$signed( -{ 1'b0,x355 } )+$signed( { 2'b0,x114 } <<<3'd1 )+$signed( -{ 1'b0,x370 } )+$signed( -{ 1'b0,x626 } )+$signed( { 2'b0,x115 } <<<3'd1 )+$signed( -{ 1'b0,x371 } )+$signed( -{ 2'b0,x627 }<<<3'd1 )+$signed(11'd40);
assign y217=temp_y[217][11] ==1'b1 ? 5'd0 :  
        temp_y[217][8] ==1'b1 ? 5'd31 : 
        temp_y[217][2]==1'b1 ? temp_y[217][7:3]+1'b1 : temp_y[217][7:3];
assign temp_y[281] = 
+$signed( -{ 1'b0,x98 } )+$signed( { 2'b0,x354 } <<<3'd1 )+$signed( -{ 1'b0,x610 } )+$signed( -{ 1'b0,x99 } )+$signed( { 2'b0,x355 } <<<3'd1 )+$signed( -{ 2'b0,x611 }<<<3'd1 )+$signed( -{ 1'b0,x114 } )+$signed( { 2'b0,x370 } <<<3'd1 )+$signed( -{ 1'b0,x626 } )+$signed( -{ 2'b0,x115 }<<<3'd1 )+$signed( { 3'b0,x371 }<<<3'd2 )+$signed( -{ 2'b0,x627 }<<<3'd1 )+$signed(11'd32);
assign y281=temp_y[281][11] ==1'b1 ? 5'd0 :  
        temp_y[281][8] ==1'b1 ? 5'd31 : 
        temp_y[281][2]==1'b1 ? temp_y[281][7:3]+1'b1 : temp_y[281][7:3];
assign temp_y[345] = 
+$signed( -{ 1'b0,x98 } )+$signed( -{ 2'b0,x354 }<<<3'd1 )+$signed( -{ 1'b0,x610 } )+$signed( { 1'b0,x99 }  )+$signed( { 2'b0,x355 } <<<3'd1 )+$signed( { 1'b0,x611 }  )+$signed( { 1'b0,x114 }  )+$signed( { 2'b0,x370 } <<<3'd1 )+$signed( { 2'b0,x626 } <<<3'd1 )+$signed( -{ 1'b0,x115 } )+$signed( -{ 2'b0,x371 }<<<3'd1 )+$signed( -{ 1'b0,x627 } )-$signed(11'd68);
assign y345=temp_y[345][11] ==1'b1 ? 5'd0 :  
        temp_y[345][8] ==1'b1 ? 5'd31 : 
        temp_y[345][2]==1'b1 ? temp_y[345][7:3]+1'b1 : temp_y[345][7:3];
assign temp_y[409] = 
+$signed( { 1'b0,x354 }  )+$signed( { 1'b0,x611 }  )+$signed( { 1'b0,x627 }  )-$signed(11'd108);
assign y409=temp_y[409][11] ==1'b1 ? 5'd0 :  
        temp_y[409][8] ==1'b1 ? 5'd31 : 
        temp_y[409][2]==1'b1 ? temp_y[409][7:3]+1'b1 : temp_y[409][7:3];
assign temp_y[473] = 
+$signed( -{ 2'b0,x98 }<<<3'd1 )+$signed( { 2'b0,x610 } <<<3'd1 )+$signed( -{ 2'b0,x99 }<<<3'd1 )+$signed( { 1'b0,x355 }  )+$signed( { 1'b0,x611 }  )+$signed( -{ 2'b0,x114 }<<<3'd1 )+$signed( { 1'b0,x370 }  )+$signed( { 1'b0,x626 }  )+$signed( -{ 1'b0,x115 } )+$signed(11'd64);
assign y473=temp_y[473][11] ==1'b1 ? 5'd0 :  
        temp_y[473][8] ==1'b1 ? 5'd31 : 
        temp_y[473][2]==1'b1 ? temp_y[473][7:3]+1'b1 : temp_y[473][7:3];
assign temp_y[537] = 
+$signed( -{ 2'b0,x98 }<<<3'd1 )+$signed( -{ 1'b0,x354 } )+$signed( -{ 3'b0,x99 }<<<3'd2)+$signed( { 1'b0,x114 }  )+$signed( { 1'b0,x370 }  )+$signed( { 3'b0,x115 }<<<3'd2 )+$signed(11'd16);
assign y537=temp_y[537][11] ==1'b1 ? 5'd0 :  
        temp_y[537][8] ==1'b1 ? 5'd31 : 
        temp_y[537][2]==1'b1 ? temp_y[537][7:3]+1'b1 : temp_y[537][7:3];
assign temp_y[601] = 
+$signed( { 2'b0,x354 } <<<3'd1 )+$signed( { 2'b0,x610 } <<<3'd1 )+$signed( -{ 1'b0,x99 } )+$signed( -{ 2'b0,x355 }<<<3'd1 )+$signed( -{ 2'b0,x611 }<<<3'd1 )+$signed( { 2'b0,x370 } <<<3'd1 )+$signed( { 1'b0,x626 }  )+$signed( -{ 2'b0,x371 }<<<3'd1 )-$signed(11'd8);
assign y601=temp_y[601][11] ==1'b1 ? 5'd0 :  
        temp_y[601][8] ==1'b1 ? 5'd31 : 
        temp_y[601][2]==1'b1 ? temp_y[601][7:3]+1'b1 : temp_y[601][7:3];
assign temp_y[26] = 
+$signed( -{ 2'b0,x356 }<<<3'd1 )+$signed( -{ 1'b0,x612 } )+$signed( { 1'b0,x101 }  )+$signed( { 1'b0,x357 }  )+$signed( { 1'b0,x613 }  )+$signed( -{ 2'b0,x372 }<<<3'd1 )+$signed( -{ 2'b0,x628 }<<<3'd1 )+$signed( { 2'b0,x373 } <<<3'd1 )+$signed( { 2'b0,x629 } <<<3'd1 )-$signed(11'd16);
assign y26=temp_y[26][11] ==1'b1 ? 5'd0 :  
        temp_y[26][8] ==1'b1 ? 5'd31 : 
        temp_y[26][2]==1'b1 ? temp_y[26][7:3]+1'b1 : temp_y[26][7:3];
assign temp_y[90] = 
+$signed( { 3'b0,x100 }<<<3'd2 )+$signed( -{ 2'b0,x356 }<<<3'd1 )+$signed( -{ 2'b0,x612 }<<<3'd1 )+$signed( { 2'b0,x101 } <<<3'd1 )+$signed( -{ 3'b0,x357 }<<<3'd2)+$signed( { 1'b0,x613 }  )+$signed( -{ 1'b0,x116 } )+$signed( { 1'b0,x628 }  )+$signed( -{ 2'b0,x117 }<<<3'd1 )+$signed( -{ 1'b0,x373 } )+$signed( { 2'b0,x629 } <<<3'd1 )+$signed(11'd24);
assign y90=temp_y[90][11] ==1'b1 ? 5'd0 :  
        temp_y[90][8] ==1'b1 ? 5'd31 : 
        temp_y[90][2]==1'b1 ? temp_y[90][7:3]+1'b1 : temp_y[90][7:3];
assign temp_y[154] = 
+$signed( { 2'b0,x100 } <<<3'd1 )+$signed( { 2'b0,x356 } <<<3'd1 )+$signed( { 1'b0,x612 }  )+$signed( { 2'b0,x101 } <<<3'd1 )+$signed( -{ 1'b0,x357 } )+$signed( { 1'b0,x613 }  )+$signed( -{ 2'b0,x116 }<<<3'd1 )+$signed( -{ 2'b0,x372 }<<<3'd1 )+$signed( -{ 1'b0,x628 } )+$signed( -{ 1'b0,x117 } )+$signed( -{ 1'b0,x373 } )+$signed( -{ 1'b0,x629 } )+$signed(11'd16);
assign y154=temp_y[154][11] ==1'b1 ? 5'd0 :  
        temp_y[154][8] ==1'b1 ? 5'd31 : 
        temp_y[154][2]==1'b1 ? temp_y[154][7:3]+1'b1 : temp_y[154][7:3];
assign temp_y[218] = 
+$signed( { 1'b0,x100 }  )+$signed( -{ 1'b0,x356 } )+$signed( { 1'b0,x101 }  )+$signed( -{ 1'b0,x357 } )+$signed( { 2'b0,x116 } <<<3'd1 )+$signed( -{ 1'b0,x372 } )+$signed( -{ 1'b0,x628 } )+$signed( { 2'b0,x117 } <<<3'd1 )+$signed( -{ 1'b0,x373 } )+$signed( -{ 2'b0,x629 }<<<3'd1 )+$signed(11'd40);
assign y218=temp_y[218][11] ==1'b1 ? 5'd0 :  
        temp_y[218][8] ==1'b1 ? 5'd31 : 
        temp_y[218][2]==1'b1 ? temp_y[218][7:3]+1'b1 : temp_y[218][7:3];
assign temp_y[282] = 
+$signed( -{ 1'b0,x100 } )+$signed( { 2'b0,x356 } <<<3'd1 )+$signed( -{ 1'b0,x612 } )+$signed( -{ 1'b0,x101 } )+$signed( { 2'b0,x357 } <<<3'd1 )+$signed( -{ 2'b0,x613 }<<<3'd1 )+$signed( -{ 1'b0,x116 } )+$signed( { 2'b0,x372 } <<<3'd1 )+$signed( -{ 1'b0,x628 } )+$signed( -{ 2'b0,x117 }<<<3'd1 )+$signed( { 3'b0,x373 }<<<3'd2 )+$signed( -{ 2'b0,x629 }<<<3'd1 )+$signed(11'd32);
assign y282=temp_y[282][11] ==1'b1 ? 5'd0 :  
        temp_y[282][8] ==1'b1 ? 5'd31 : 
        temp_y[282][2]==1'b1 ? temp_y[282][7:3]+1'b1 : temp_y[282][7:3];
assign temp_y[346] = 
+$signed( -{ 1'b0,x100 } )+$signed( -{ 2'b0,x356 }<<<3'd1 )+$signed( -{ 1'b0,x612 } )+$signed( { 1'b0,x101 }  )+$signed( { 2'b0,x357 } <<<3'd1 )+$signed( { 1'b0,x613 }  )+$signed( { 1'b0,x116 }  )+$signed( { 2'b0,x372 } <<<3'd1 )+$signed( { 2'b0,x628 } <<<3'd1 )+$signed( -{ 1'b0,x117 } )+$signed( -{ 2'b0,x373 }<<<3'd1 )+$signed( -{ 1'b0,x629 } )-$signed(11'd68);
assign y346=temp_y[346][11] ==1'b1 ? 5'd0 :  
        temp_y[346][8] ==1'b1 ? 5'd31 : 
        temp_y[346][2]==1'b1 ? temp_y[346][7:3]+1'b1 : temp_y[346][7:3];
assign temp_y[410] = 
+$signed( { 1'b0,x356 }  )+$signed( { 1'b0,x613 }  )+$signed( { 1'b0,x629 }  )-$signed(11'd108);
assign y410=temp_y[410][11] ==1'b1 ? 5'd0 :  
        temp_y[410][8] ==1'b1 ? 5'd31 : 
        temp_y[410][2]==1'b1 ? temp_y[410][7:3]+1'b1 : temp_y[410][7:3];
assign temp_y[474] = 
+$signed( -{ 2'b0,x100 }<<<3'd1 )+$signed( { 2'b0,x612 } <<<3'd1 )+$signed( -{ 2'b0,x101 }<<<3'd1 )+$signed( { 1'b0,x357 }  )+$signed( { 1'b0,x613 }  )+$signed( -{ 2'b0,x116 }<<<3'd1 )+$signed( { 1'b0,x372 }  )+$signed( { 1'b0,x628 }  )+$signed( -{ 1'b0,x117 } )+$signed(11'd64);
assign y474=temp_y[474][11] ==1'b1 ? 5'd0 :  
        temp_y[474][8] ==1'b1 ? 5'd31 : 
        temp_y[474][2]==1'b1 ? temp_y[474][7:3]+1'b1 : temp_y[474][7:3];
assign temp_y[538] = 
+$signed( -{ 2'b0,x100 }<<<3'd1 )+$signed( -{ 1'b0,x356 } )+$signed( -{ 3'b0,x101 }<<<3'd2)+$signed( { 1'b0,x116 }  )+$signed( { 1'b0,x372 }  )+$signed( { 3'b0,x117 }<<<3'd2 )+$signed(11'd16);
assign y538=temp_y[538][11] ==1'b1 ? 5'd0 :  
        temp_y[538][8] ==1'b1 ? 5'd31 : 
        temp_y[538][2]==1'b1 ? temp_y[538][7:3]+1'b1 : temp_y[538][7:3];
assign temp_y[602] = 
+$signed( { 2'b0,x356 } <<<3'd1 )+$signed( { 2'b0,x612 } <<<3'd1 )+$signed( -{ 1'b0,x101 } )+$signed( -{ 2'b0,x357 }<<<3'd1 )+$signed( -{ 2'b0,x613 }<<<3'd1 )+$signed( { 2'b0,x372 } <<<3'd1 )+$signed( { 1'b0,x628 }  )+$signed( -{ 2'b0,x373 }<<<3'd1 )-$signed(11'd8);
assign y602=temp_y[602][11] ==1'b1 ? 5'd0 :  
        temp_y[602][8] ==1'b1 ? 5'd31 : 
        temp_y[602][2]==1'b1 ? temp_y[602][7:3]+1'b1 : temp_y[602][7:3];
assign temp_y[27] = 
+$signed( -{ 2'b0,x358 }<<<3'd1 )+$signed( -{ 1'b0,x614 } )+$signed( { 1'b0,x103 }  )+$signed( { 1'b0,x359 }  )+$signed( { 1'b0,x615 }  )+$signed( -{ 2'b0,x374 }<<<3'd1 )+$signed( -{ 2'b0,x630 }<<<3'd1 )+$signed( { 2'b0,x375 } <<<3'd1 )+$signed( { 2'b0,x631 } <<<3'd1 )-$signed(11'd16);
assign y27=temp_y[27][11] ==1'b1 ? 5'd0 :  
        temp_y[27][8] ==1'b1 ? 5'd31 : 
        temp_y[27][2]==1'b1 ? temp_y[27][7:3]+1'b1 : temp_y[27][7:3];
assign temp_y[91] = 
+$signed( { 3'b0,x102 }<<<3'd2 )+$signed( -{ 2'b0,x358 }<<<3'd1 )+$signed( -{ 2'b0,x614 }<<<3'd1 )+$signed( { 2'b0,x103 } <<<3'd1 )+$signed( -{ 3'b0,x359 }<<<3'd2)+$signed( { 1'b0,x615 }  )+$signed( -{ 1'b0,x118 } )+$signed( { 1'b0,x630 }  )+$signed( -{ 2'b0,x119 }<<<3'd1 )+$signed( -{ 1'b0,x375 } )+$signed( { 2'b0,x631 } <<<3'd1 )+$signed(11'd24);
assign y91=temp_y[91][11] ==1'b1 ? 5'd0 :  
        temp_y[91][8] ==1'b1 ? 5'd31 : 
        temp_y[91][2]==1'b1 ? temp_y[91][7:3]+1'b1 : temp_y[91][7:3];
assign temp_y[155] = 
+$signed( { 2'b0,x102 } <<<3'd1 )+$signed( { 2'b0,x358 } <<<3'd1 )+$signed( { 1'b0,x614 }  )+$signed( { 2'b0,x103 } <<<3'd1 )+$signed( -{ 1'b0,x359 } )+$signed( { 1'b0,x615 }  )+$signed( -{ 2'b0,x118 }<<<3'd1 )+$signed( -{ 2'b0,x374 }<<<3'd1 )+$signed( -{ 1'b0,x630 } )+$signed( -{ 1'b0,x119 } )+$signed( -{ 1'b0,x375 } )+$signed( -{ 1'b0,x631 } )+$signed(11'd16);
assign y155=temp_y[155][11] ==1'b1 ? 5'd0 :  
        temp_y[155][8] ==1'b1 ? 5'd31 : 
        temp_y[155][2]==1'b1 ? temp_y[155][7:3]+1'b1 : temp_y[155][7:3];
assign temp_y[219] = 
+$signed( { 1'b0,x102 }  )+$signed( -{ 1'b0,x358 } )+$signed( { 1'b0,x103 }  )+$signed( -{ 1'b0,x359 } )+$signed( { 2'b0,x118 } <<<3'd1 )+$signed( -{ 1'b0,x374 } )+$signed( -{ 1'b0,x630 } )+$signed( { 2'b0,x119 } <<<3'd1 )+$signed( -{ 1'b0,x375 } )+$signed( -{ 2'b0,x631 }<<<3'd1 )+$signed(11'd40);
assign y219=temp_y[219][11] ==1'b1 ? 5'd0 :  
        temp_y[219][8] ==1'b1 ? 5'd31 : 
        temp_y[219][2]==1'b1 ? temp_y[219][7:3]+1'b1 : temp_y[219][7:3];
assign temp_y[283] = 
+$signed( -{ 1'b0,x102 } )+$signed( { 2'b0,x358 } <<<3'd1 )+$signed( -{ 1'b0,x614 } )+$signed( -{ 1'b0,x103 } )+$signed( { 2'b0,x359 } <<<3'd1 )+$signed( -{ 2'b0,x615 }<<<3'd1 )+$signed( -{ 1'b0,x118 } )+$signed( { 2'b0,x374 } <<<3'd1 )+$signed( -{ 1'b0,x630 } )+$signed( -{ 2'b0,x119 }<<<3'd1 )+$signed( { 3'b0,x375 }<<<3'd2 )+$signed( -{ 2'b0,x631 }<<<3'd1 )+$signed(11'd32);
assign y283=temp_y[283][11] ==1'b1 ? 5'd0 :  
        temp_y[283][8] ==1'b1 ? 5'd31 : 
        temp_y[283][2]==1'b1 ? temp_y[283][7:3]+1'b1 : temp_y[283][7:3];
assign temp_y[347] = 
+$signed( -{ 1'b0,x102 } )+$signed( -{ 2'b0,x358 }<<<3'd1 )+$signed( -{ 1'b0,x614 } )+$signed( { 1'b0,x103 }  )+$signed( { 2'b0,x359 } <<<3'd1 )+$signed( { 1'b0,x615 }  )+$signed( { 1'b0,x118 }  )+$signed( { 2'b0,x374 } <<<3'd1 )+$signed( { 2'b0,x630 } <<<3'd1 )+$signed( -{ 1'b0,x119 } )+$signed( -{ 2'b0,x375 }<<<3'd1 )+$signed( -{ 1'b0,x631 } )-$signed(11'd68);
assign y347=temp_y[347][11] ==1'b1 ? 5'd0 :  
        temp_y[347][8] ==1'b1 ? 5'd31 : 
        temp_y[347][2]==1'b1 ? temp_y[347][7:3]+1'b1 : temp_y[347][7:3];
assign temp_y[411] = 
+$signed( { 1'b0,x358 }  )+$signed( { 1'b0,x615 }  )+$signed( { 1'b0,x631 }  )-$signed(11'd108);
assign y411=temp_y[411][11] ==1'b1 ? 5'd0 :  
        temp_y[411][8] ==1'b1 ? 5'd31 : 
        temp_y[411][2]==1'b1 ? temp_y[411][7:3]+1'b1 : temp_y[411][7:3];
assign temp_y[475] = 
+$signed( -{ 2'b0,x102 }<<<3'd1 )+$signed( { 2'b0,x614 } <<<3'd1 )+$signed( -{ 2'b0,x103 }<<<3'd1 )+$signed( { 1'b0,x359 }  )+$signed( { 1'b0,x615 }  )+$signed( -{ 2'b0,x118 }<<<3'd1 )+$signed( { 1'b0,x374 }  )+$signed( { 1'b0,x630 }  )+$signed( -{ 1'b0,x119 } )+$signed(11'd64);
assign y475=temp_y[475][11] ==1'b1 ? 5'd0 :  
        temp_y[475][8] ==1'b1 ? 5'd31 : 
        temp_y[475][2]==1'b1 ? temp_y[475][7:3]+1'b1 : temp_y[475][7:3];
assign temp_y[539] = 
+$signed( -{ 2'b0,x102 }<<<3'd1 )+$signed( -{ 1'b0,x358 } )+$signed( -{ 3'b0,x103 }<<<3'd2)+$signed( { 1'b0,x118 }  )+$signed( { 1'b0,x374 }  )+$signed( { 3'b0,x119 }<<<3'd2 )+$signed(11'd16);
assign y539=temp_y[539][11] ==1'b1 ? 5'd0 :  
        temp_y[539][8] ==1'b1 ? 5'd31 : 
        temp_y[539][2]==1'b1 ? temp_y[539][7:3]+1'b1 : temp_y[539][7:3];
assign temp_y[603] = 
+$signed( { 2'b0,x358 } <<<3'd1 )+$signed( { 2'b0,x614 } <<<3'd1 )+$signed( -{ 1'b0,x103 } )+$signed( -{ 2'b0,x359 }<<<3'd1 )+$signed( -{ 2'b0,x615 }<<<3'd1 )+$signed( { 2'b0,x374 } <<<3'd1 )+$signed( { 1'b0,x630 }  )+$signed( -{ 2'b0,x375 }<<<3'd1 )-$signed(11'd8);
assign y603=temp_y[603][11] ==1'b1 ? 5'd0 :  
        temp_y[603][8] ==1'b1 ? 5'd31 : 
        temp_y[603][2]==1'b1 ? temp_y[603][7:3]+1'b1 : temp_y[603][7:3];
assign temp_y[28] = 
+$signed( -{ 2'b0,x360 }<<<3'd1 )+$signed( -{ 1'b0,x616 } )+$signed( { 1'b0,x105 }  )+$signed( { 1'b0,x361 }  )+$signed( { 1'b0,x617 }  )+$signed( -{ 2'b0,x376 }<<<3'd1 )+$signed( -{ 2'b0,x632 }<<<3'd1 )+$signed( { 2'b0,x377 } <<<3'd1 )+$signed( { 2'b0,x633 } <<<3'd1 )-$signed(11'd16);
assign y28=temp_y[28][11] ==1'b1 ? 5'd0 :  
        temp_y[28][8] ==1'b1 ? 5'd31 : 
        temp_y[28][2]==1'b1 ? temp_y[28][7:3]+1'b1 : temp_y[28][7:3];
assign temp_y[92] = 
+$signed( { 3'b0,x104 }<<<3'd2 )+$signed( -{ 2'b0,x360 }<<<3'd1 )+$signed( -{ 2'b0,x616 }<<<3'd1 )+$signed( { 2'b0,x105 } <<<3'd1 )+$signed( -{ 3'b0,x361 }<<<3'd2)+$signed( { 1'b0,x617 }  )+$signed( -{ 1'b0,x120 } )+$signed( { 1'b0,x632 }  )+$signed( -{ 2'b0,x121 }<<<3'd1 )+$signed( -{ 1'b0,x377 } )+$signed( { 2'b0,x633 } <<<3'd1 )+$signed(11'd24);
assign y92=temp_y[92][11] ==1'b1 ? 5'd0 :  
        temp_y[92][8] ==1'b1 ? 5'd31 : 
        temp_y[92][2]==1'b1 ? temp_y[92][7:3]+1'b1 : temp_y[92][7:3];
assign temp_y[156] = 
+$signed( { 2'b0,x104 } <<<3'd1 )+$signed( { 2'b0,x360 } <<<3'd1 )+$signed( { 1'b0,x616 }  )+$signed( { 2'b0,x105 } <<<3'd1 )+$signed( -{ 1'b0,x361 } )+$signed( { 1'b0,x617 }  )+$signed( -{ 2'b0,x120 }<<<3'd1 )+$signed( -{ 2'b0,x376 }<<<3'd1 )+$signed( -{ 1'b0,x632 } )+$signed( -{ 1'b0,x121 } )+$signed( -{ 1'b0,x377 } )+$signed( -{ 1'b0,x633 } )+$signed(11'd16);
assign y156=temp_y[156][11] ==1'b1 ? 5'd0 :  
        temp_y[156][8] ==1'b1 ? 5'd31 : 
        temp_y[156][2]==1'b1 ? temp_y[156][7:3]+1'b1 : temp_y[156][7:3];
assign temp_y[220] = 
+$signed( { 1'b0,x104 }  )+$signed( -{ 1'b0,x360 } )+$signed( { 1'b0,x105 }  )+$signed( -{ 1'b0,x361 } )+$signed( { 2'b0,x120 } <<<3'd1 )+$signed( -{ 1'b0,x376 } )+$signed( -{ 1'b0,x632 } )+$signed( { 2'b0,x121 } <<<3'd1 )+$signed( -{ 1'b0,x377 } )+$signed( -{ 2'b0,x633 }<<<3'd1 )+$signed(11'd40);
assign y220=temp_y[220][11] ==1'b1 ? 5'd0 :  
        temp_y[220][8] ==1'b1 ? 5'd31 : 
        temp_y[220][2]==1'b1 ? temp_y[220][7:3]+1'b1 : temp_y[220][7:3];
assign temp_y[284] = 
+$signed( -{ 1'b0,x104 } )+$signed( { 2'b0,x360 } <<<3'd1 )+$signed( -{ 1'b0,x616 } )+$signed( -{ 1'b0,x105 } )+$signed( { 2'b0,x361 } <<<3'd1 )+$signed( -{ 2'b0,x617 }<<<3'd1 )+$signed( -{ 1'b0,x120 } )+$signed( { 2'b0,x376 } <<<3'd1 )+$signed( -{ 1'b0,x632 } )+$signed( -{ 2'b0,x121 }<<<3'd1 )+$signed( { 3'b0,x377 }<<<3'd2 )+$signed( -{ 2'b0,x633 }<<<3'd1 )+$signed(11'd32);
assign y284=temp_y[284][11] ==1'b1 ? 5'd0 :  
        temp_y[284][8] ==1'b1 ? 5'd31 : 
        temp_y[284][2]==1'b1 ? temp_y[284][7:3]+1'b1 : temp_y[284][7:3];
assign temp_y[348] = 
+$signed( -{ 1'b0,x104 } )+$signed( -{ 2'b0,x360 }<<<3'd1 )+$signed( -{ 1'b0,x616 } )+$signed( { 1'b0,x105 }  )+$signed( { 2'b0,x361 } <<<3'd1 )+$signed( { 1'b0,x617 }  )+$signed( { 1'b0,x120 }  )+$signed( { 2'b0,x376 } <<<3'd1 )+$signed( { 2'b0,x632 } <<<3'd1 )+$signed( -{ 1'b0,x121 } )+$signed( -{ 2'b0,x377 }<<<3'd1 )+$signed( -{ 1'b0,x633 } )-$signed(11'd68);
assign y348=temp_y[348][11] ==1'b1 ? 5'd0 :  
        temp_y[348][8] ==1'b1 ? 5'd31 : 
        temp_y[348][2]==1'b1 ? temp_y[348][7:3]+1'b1 : temp_y[348][7:3];
assign temp_y[412] = 
+$signed( { 1'b0,x360 }  )+$signed( { 1'b0,x617 }  )+$signed( { 1'b0,x633 }  )-$signed(11'd108);
assign y412=temp_y[412][11] ==1'b1 ? 5'd0 :  
        temp_y[412][8] ==1'b1 ? 5'd31 : 
        temp_y[412][2]==1'b1 ? temp_y[412][7:3]+1'b1 : temp_y[412][7:3];
assign temp_y[476] = 
+$signed( -{ 2'b0,x104 }<<<3'd1 )+$signed( { 2'b0,x616 } <<<3'd1 )+$signed( -{ 2'b0,x105 }<<<3'd1 )+$signed( { 1'b0,x361 }  )+$signed( { 1'b0,x617 }  )+$signed( -{ 2'b0,x120 }<<<3'd1 )+$signed( { 1'b0,x376 }  )+$signed( { 1'b0,x632 }  )+$signed( -{ 1'b0,x121 } )+$signed(11'd64);
assign y476=temp_y[476][11] ==1'b1 ? 5'd0 :  
        temp_y[476][8] ==1'b1 ? 5'd31 : 
        temp_y[476][2]==1'b1 ? temp_y[476][7:3]+1'b1 : temp_y[476][7:3];
assign temp_y[540] = 
+$signed( -{ 2'b0,x104 }<<<3'd1 )+$signed( -{ 1'b0,x360 } )+$signed( -{ 3'b0,x105 }<<<3'd2)+$signed( { 1'b0,x120 }  )+$signed( { 1'b0,x376 }  )+$signed( { 3'b0,x121 }<<<3'd2 )+$signed(11'd16);
assign y540=temp_y[540][11] ==1'b1 ? 5'd0 :  
        temp_y[540][8] ==1'b1 ? 5'd31 : 
        temp_y[540][2]==1'b1 ? temp_y[540][7:3]+1'b1 : temp_y[540][7:3];
assign temp_y[604] = 
+$signed( { 2'b0,x360 } <<<3'd1 )+$signed( { 2'b0,x616 } <<<3'd1 )+$signed( -{ 1'b0,x105 } )+$signed( -{ 2'b0,x361 }<<<3'd1 )+$signed( -{ 2'b0,x617 }<<<3'd1 )+$signed( { 2'b0,x376 } <<<3'd1 )+$signed( { 1'b0,x632 }  )+$signed( -{ 2'b0,x377 }<<<3'd1 )-$signed(11'd8);
assign y604=temp_y[604][11] ==1'b1 ? 5'd0 :  
        temp_y[604][8] ==1'b1 ? 5'd31 : 
        temp_y[604][2]==1'b1 ? temp_y[604][7:3]+1'b1 : temp_y[604][7:3];
assign temp_y[29] = 
+$signed( -{ 2'b0,x362 }<<<3'd1 )+$signed( -{ 1'b0,x618 } )+$signed( { 1'b0,x107 }  )+$signed( { 1'b0,x363 }  )+$signed( { 1'b0,x619 }  )+$signed( -{ 2'b0,x378 }<<<3'd1 )+$signed( -{ 2'b0,x634 }<<<3'd1 )+$signed( { 2'b0,x379 } <<<3'd1 )+$signed( { 2'b0,x635 } <<<3'd1 )-$signed(11'd16);
assign y29=temp_y[29][11] ==1'b1 ? 5'd0 :  
        temp_y[29][8] ==1'b1 ? 5'd31 : 
        temp_y[29][2]==1'b1 ? temp_y[29][7:3]+1'b1 : temp_y[29][7:3];
assign temp_y[93] = 
+$signed( { 3'b0,x106 }<<<3'd2 )+$signed( -{ 2'b0,x362 }<<<3'd1 )+$signed( -{ 2'b0,x618 }<<<3'd1 )+$signed( { 2'b0,x107 } <<<3'd1 )+$signed( -{ 3'b0,x363 }<<<3'd2)+$signed( { 1'b0,x619 }  )+$signed( -{ 1'b0,x122 } )+$signed( { 1'b0,x634 }  )+$signed( -{ 2'b0,x123 }<<<3'd1 )+$signed( -{ 1'b0,x379 } )+$signed( { 2'b0,x635 } <<<3'd1 )+$signed(11'd24);
assign y93=temp_y[93][11] ==1'b1 ? 5'd0 :  
        temp_y[93][8] ==1'b1 ? 5'd31 : 
        temp_y[93][2]==1'b1 ? temp_y[93][7:3]+1'b1 : temp_y[93][7:3];
assign temp_y[157] = 
+$signed( { 2'b0,x106 } <<<3'd1 )+$signed( { 2'b0,x362 } <<<3'd1 )+$signed( { 1'b0,x618 }  )+$signed( { 2'b0,x107 } <<<3'd1 )+$signed( -{ 1'b0,x363 } )+$signed( { 1'b0,x619 }  )+$signed( -{ 2'b0,x122 }<<<3'd1 )+$signed( -{ 2'b0,x378 }<<<3'd1 )+$signed( -{ 1'b0,x634 } )+$signed( -{ 1'b0,x123 } )+$signed( -{ 1'b0,x379 } )+$signed( -{ 1'b0,x635 } )+$signed(11'd16);
assign y157=temp_y[157][11] ==1'b1 ? 5'd0 :  
        temp_y[157][8] ==1'b1 ? 5'd31 : 
        temp_y[157][2]==1'b1 ? temp_y[157][7:3]+1'b1 : temp_y[157][7:3];
assign temp_y[221] = 
+$signed( { 1'b0,x106 }  )+$signed( -{ 1'b0,x362 } )+$signed( { 1'b0,x107 }  )+$signed( -{ 1'b0,x363 } )+$signed( { 2'b0,x122 } <<<3'd1 )+$signed( -{ 1'b0,x378 } )+$signed( -{ 1'b0,x634 } )+$signed( { 2'b0,x123 } <<<3'd1 )+$signed( -{ 1'b0,x379 } )+$signed( -{ 2'b0,x635 }<<<3'd1 )+$signed(11'd40);
assign y221=temp_y[221][11] ==1'b1 ? 5'd0 :  
        temp_y[221][8] ==1'b1 ? 5'd31 : 
        temp_y[221][2]==1'b1 ? temp_y[221][7:3]+1'b1 : temp_y[221][7:3];
assign temp_y[285] = 
+$signed( -{ 1'b0,x106 } )+$signed( { 2'b0,x362 } <<<3'd1 )+$signed( -{ 1'b0,x618 } )+$signed( -{ 1'b0,x107 } )+$signed( { 2'b0,x363 } <<<3'd1 )+$signed( -{ 2'b0,x619 }<<<3'd1 )+$signed( -{ 1'b0,x122 } )+$signed( { 2'b0,x378 } <<<3'd1 )+$signed( -{ 1'b0,x634 } )+$signed( -{ 2'b0,x123 }<<<3'd1 )+$signed( { 3'b0,x379 }<<<3'd2 )+$signed( -{ 2'b0,x635 }<<<3'd1 )+$signed(11'd32);
assign y285=temp_y[285][11] ==1'b1 ? 5'd0 :  
        temp_y[285][8] ==1'b1 ? 5'd31 : 
        temp_y[285][2]==1'b1 ? temp_y[285][7:3]+1'b1 : temp_y[285][7:3];
assign temp_y[349] = 
+$signed( -{ 1'b0,x106 } )+$signed( -{ 2'b0,x362 }<<<3'd1 )+$signed( -{ 1'b0,x618 } )+$signed( { 1'b0,x107 }  )+$signed( { 2'b0,x363 } <<<3'd1 )+$signed( { 1'b0,x619 }  )+$signed( { 1'b0,x122 }  )+$signed( { 2'b0,x378 } <<<3'd1 )+$signed( { 2'b0,x634 } <<<3'd1 )+$signed( -{ 1'b0,x123 } )+$signed( -{ 2'b0,x379 }<<<3'd1 )+$signed( -{ 1'b0,x635 } )-$signed(11'd68);
assign y349=temp_y[349][11] ==1'b1 ? 5'd0 :  
        temp_y[349][8] ==1'b1 ? 5'd31 : 
        temp_y[349][2]==1'b1 ? temp_y[349][7:3]+1'b1 : temp_y[349][7:3];
assign temp_y[413] = 
+$signed( { 1'b0,x362 }  )+$signed( { 1'b0,x619 }  )+$signed( { 1'b0,x635 }  )-$signed(11'd108);
assign y413=temp_y[413][11] ==1'b1 ? 5'd0 :  
        temp_y[413][8] ==1'b1 ? 5'd31 : 
        temp_y[413][2]==1'b1 ? temp_y[413][7:3]+1'b1 : temp_y[413][7:3];
assign temp_y[477] = 
+$signed( -{ 2'b0,x106 }<<<3'd1 )+$signed( { 2'b0,x618 } <<<3'd1 )+$signed( -{ 2'b0,x107 }<<<3'd1 )+$signed( { 1'b0,x363 }  )+$signed( { 1'b0,x619 }  )+$signed( -{ 2'b0,x122 }<<<3'd1 )+$signed( { 1'b0,x378 }  )+$signed( { 1'b0,x634 }  )+$signed( -{ 1'b0,x123 } )+$signed(11'd64);
assign y477=temp_y[477][11] ==1'b1 ? 5'd0 :  
        temp_y[477][8] ==1'b1 ? 5'd31 : 
        temp_y[477][2]==1'b1 ? temp_y[477][7:3]+1'b1 : temp_y[477][7:3];
assign temp_y[541] = 
+$signed( -{ 2'b0,x106 }<<<3'd1 )+$signed( -{ 1'b0,x362 } )+$signed( -{ 3'b0,x107 }<<<3'd2)+$signed( { 1'b0,x122 }  )+$signed( { 1'b0,x378 }  )+$signed( { 3'b0,x123 }<<<3'd2 )+$signed(11'd16);
assign y541=temp_y[541][11] ==1'b1 ? 5'd0 :  
        temp_y[541][8] ==1'b1 ? 5'd31 : 
        temp_y[541][2]==1'b1 ? temp_y[541][7:3]+1'b1 : temp_y[541][7:3];
assign temp_y[605] = 
+$signed( { 2'b0,x362 } <<<3'd1 )+$signed( { 2'b0,x618 } <<<3'd1 )+$signed( -{ 1'b0,x107 } )+$signed( -{ 2'b0,x363 }<<<3'd1 )+$signed( -{ 2'b0,x619 }<<<3'd1 )+$signed( { 2'b0,x378 } <<<3'd1 )+$signed( { 1'b0,x634 }  )+$signed( -{ 2'b0,x379 }<<<3'd1 )-$signed(11'd8);
assign y605=temp_y[605][11] ==1'b1 ? 5'd0 :  
        temp_y[605][8] ==1'b1 ? 5'd31 : 
        temp_y[605][2]==1'b1 ? temp_y[605][7:3]+1'b1 : temp_y[605][7:3];
assign temp_y[30] = 
+$signed( -{ 2'b0,x364 }<<<3'd1 )+$signed( -{ 1'b0,x620 } )+$signed( { 1'b0,x109 }  )+$signed( { 1'b0,x365 }  )+$signed( { 1'b0,x621 }  )+$signed( -{ 2'b0,x380 }<<<3'd1 )+$signed( -{ 2'b0,x636 }<<<3'd1 )+$signed( { 2'b0,x381 } <<<3'd1 )+$signed( { 2'b0,x637 } <<<3'd1 )-$signed(11'd16);
assign y30=temp_y[30][11] ==1'b1 ? 5'd0 :  
        temp_y[30][8] ==1'b1 ? 5'd31 : 
        temp_y[30][2]==1'b1 ? temp_y[30][7:3]+1'b1 : temp_y[30][7:3];
assign temp_y[94] = 
+$signed( { 3'b0,x108 }<<<3'd2 )+$signed( -{ 2'b0,x364 }<<<3'd1 )+$signed( -{ 2'b0,x620 }<<<3'd1 )+$signed( { 2'b0,x109 } <<<3'd1 )+$signed( -{ 3'b0,x365 }<<<3'd2)+$signed( { 1'b0,x621 }  )+$signed( -{ 1'b0,x124 } )+$signed( { 1'b0,x636 }  )+$signed( -{ 2'b0,x125 }<<<3'd1 )+$signed( -{ 1'b0,x381 } )+$signed( { 2'b0,x637 } <<<3'd1 )+$signed(11'd24);
assign y94=temp_y[94][11] ==1'b1 ? 5'd0 :  
        temp_y[94][8] ==1'b1 ? 5'd31 : 
        temp_y[94][2]==1'b1 ? temp_y[94][7:3]+1'b1 : temp_y[94][7:3];
assign temp_y[158] = 
+$signed( { 2'b0,x108 } <<<3'd1 )+$signed( { 2'b0,x364 } <<<3'd1 )+$signed( { 1'b0,x620 }  )+$signed( { 2'b0,x109 } <<<3'd1 )+$signed( -{ 1'b0,x365 } )+$signed( { 1'b0,x621 }  )+$signed( -{ 2'b0,x124 }<<<3'd1 )+$signed( -{ 2'b0,x380 }<<<3'd1 )+$signed( -{ 1'b0,x636 } )+$signed( -{ 1'b0,x125 } )+$signed( -{ 1'b0,x381 } )+$signed( -{ 1'b0,x637 } )+$signed(11'd16);
assign y158=temp_y[158][11] ==1'b1 ? 5'd0 :  
        temp_y[158][8] ==1'b1 ? 5'd31 : 
        temp_y[158][2]==1'b1 ? temp_y[158][7:3]+1'b1 : temp_y[158][7:3];
assign temp_y[222] = 
+$signed( { 1'b0,x108 }  )+$signed( -{ 1'b0,x364 } )+$signed( { 1'b0,x109 }  )+$signed( -{ 1'b0,x365 } )+$signed( { 2'b0,x124 } <<<3'd1 )+$signed( -{ 1'b0,x380 } )+$signed( -{ 1'b0,x636 } )+$signed( { 2'b0,x125 } <<<3'd1 )+$signed( -{ 1'b0,x381 } )+$signed( -{ 2'b0,x637 }<<<3'd1 )+$signed(11'd40);
assign y222=temp_y[222][11] ==1'b1 ? 5'd0 :  
        temp_y[222][8] ==1'b1 ? 5'd31 : 
        temp_y[222][2]==1'b1 ? temp_y[222][7:3]+1'b1 : temp_y[222][7:3];
assign temp_y[286] = 
+$signed( -{ 1'b0,x108 } )+$signed( { 2'b0,x364 } <<<3'd1 )+$signed( -{ 1'b0,x620 } )+$signed( -{ 1'b0,x109 } )+$signed( { 2'b0,x365 } <<<3'd1 )+$signed( -{ 2'b0,x621 }<<<3'd1 )+$signed( -{ 1'b0,x124 } )+$signed( { 2'b0,x380 } <<<3'd1 )+$signed( -{ 1'b0,x636 } )+$signed( -{ 2'b0,x125 }<<<3'd1 )+$signed( { 3'b0,x381 }<<<3'd2 )+$signed( -{ 2'b0,x637 }<<<3'd1 )+$signed(11'd32);
assign y286=temp_y[286][11] ==1'b1 ? 5'd0 :  
        temp_y[286][8] ==1'b1 ? 5'd31 : 
        temp_y[286][2]==1'b1 ? temp_y[286][7:3]+1'b1 : temp_y[286][7:3];
assign temp_y[350] = 
+$signed( -{ 1'b0,x108 } )+$signed( -{ 2'b0,x364 }<<<3'd1 )+$signed( -{ 1'b0,x620 } )+$signed( { 1'b0,x109 }  )+$signed( { 2'b0,x365 } <<<3'd1 )+$signed( { 1'b0,x621 }  )+$signed( { 1'b0,x124 }  )+$signed( { 2'b0,x380 } <<<3'd1 )+$signed( { 2'b0,x636 } <<<3'd1 )+$signed( -{ 1'b0,x125 } )+$signed( -{ 2'b0,x381 }<<<3'd1 )+$signed( -{ 1'b0,x637 } )-$signed(11'd68);
assign y350=temp_y[350][11] ==1'b1 ? 5'd0 :  
        temp_y[350][8] ==1'b1 ? 5'd31 : 
        temp_y[350][2]==1'b1 ? temp_y[350][7:3]+1'b1 : temp_y[350][7:3];
assign temp_y[414] = 
+$signed( { 1'b0,x364 }  )+$signed( { 1'b0,x621 }  )+$signed( { 1'b0,x637 }  )-$signed(11'd108);
assign y414=temp_y[414][11] ==1'b1 ? 5'd0 :  
        temp_y[414][8] ==1'b1 ? 5'd31 : 
        temp_y[414][2]==1'b1 ? temp_y[414][7:3]+1'b1 : temp_y[414][7:3];
assign temp_y[478] = 
+$signed( -{ 2'b0,x108 }<<<3'd1 )+$signed( { 2'b0,x620 } <<<3'd1 )+$signed( -{ 2'b0,x109 }<<<3'd1 )+$signed( { 1'b0,x365 }  )+$signed( { 1'b0,x621 }  )+$signed( -{ 2'b0,x124 }<<<3'd1 )+$signed( { 1'b0,x380 }  )+$signed( { 1'b0,x636 }  )+$signed( -{ 1'b0,x125 } )+$signed(11'd64);
assign y478=temp_y[478][11] ==1'b1 ? 5'd0 :  
        temp_y[478][8] ==1'b1 ? 5'd31 : 
        temp_y[478][2]==1'b1 ? temp_y[478][7:3]+1'b1 : temp_y[478][7:3];
assign temp_y[542] = 
+$signed( -{ 2'b0,x108 }<<<3'd1 )+$signed( -{ 1'b0,x364 } )+$signed( -{ 3'b0,x109 }<<<3'd2)+$signed( { 1'b0,x124 }  )+$signed( { 1'b0,x380 }  )+$signed( { 3'b0,x125 }<<<3'd2 )+$signed(11'd16);
assign y542=temp_y[542][11] ==1'b1 ? 5'd0 :  
        temp_y[542][8] ==1'b1 ? 5'd31 : 
        temp_y[542][2]==1'b1 ? temp_y[542][7:3]+1'b1 : temp_y[542][7:3];
assign temp_y[606] = 
+$signed( { 2'b0,x364 } <<<3'd1 )+$signed( { 2'b0,x620 } <<<3'd1 )+$signed( -{ 1'b0,x109 } )+$signed( -{ 2'b0,x365 }<<<3'd1 )+$signed( -{ 2'b0,x621 }<<<3'd1 )+$signed( { 2'b0,x380 } <<<3'd1 )+$signed( { 1'b0,x636 }  )+$signed( -{ 2'b0,x381 }<<<3'd1 )-$signed(11'd8);
assign y606=temp_y[606][11] ==1'b1 ? 5'd0 :  
        temp_y[606][8] ==1'b1 ? 5'd31 : 
        temp_y[606][2]==1'b1 ? temp_y[606][7:3]+1'b1 : temp_y[606][7:3];
assign temp_y[31] = 
+$signed( -{ 2'b0,x366 }<<<3'd1 )+$signed( -{ 1'b0,x622 } )+$signed( { 1'b0,x111 }  )+$signed( { 1'b0,x367 }  )+$signed( { 1'b0,x623 }  )+$signed( -{ 2'b0,x382 }<<<3'd1 )+$signed( -{ 2'b0,x638 }<<<3'd1 )+$signed( { 2'b0,x383 } <<<3'd1 )+$signed( { 2'b0,x639 } <<<3'd1 )-$signed(11'd16);
assign y31=temp_y[31][11] ==1'b1 ? 5'd0 :  
        temp_y[31][8] ==1'b1 ? 5'd31 : 
        temp_y[31][2]==1'b1 ? temp_y[31][7:3]+1'b1 : temp_y[31][7:3];
assign temp_y[95] = 
+$signed( { 3'b0,x110 }<<<3'd2 )+$signed( -{ 2'b0,x366 }<<<3'd1 )+$signed( -{ 2'b0,x622 }<<<3'd1 )+$signed( { 2'b0,x111 } <<<3'd1 )+$signed( -{ 3'b0,x367 }<<<3'd2)+$signed( { 1'b0,x623 }  )+$signed( -{ 1'b0,x126 } )+$signed( { 1'b0,x638 }  )+$signed( -{ 2'b0,x127 }<<<3'd1 )+$signed( -{ 1'b0,x383 } )+$signed( { 2'b0,x639 } <<<3'd1 )+$signed(11'd24);
assign y95=temp_y[95][11] ==1'b1 ? 5'd0 :  
        temp_y[95][8] ==1'b1 ? 5'd31 : 
        temp_y[95][2]==1'b1 ? temp_y[95][7:3]+1'b1 : temp_y[95][7:3];
assign temp_y[159] = 
+$signed( { 2'b0,x110 } <<<3'd1 )+$signed( { 2'b0,x366 } <<<3'd1 )+$signed( { 1'b0,x622 }  )+$signed( { 2'b0,x111 } <<<3'd1 )+$signed( -{ 1'b0,x367 } )+$signed( { 1'b0,x623 }  )+$signed( -{ 2'b0,x126 }<<<3'd1 )+$signed( -{ 2'b0,x382 }<<<3'd1 )+$signed( -{ 1'b0,x638 } )+$signed( -{ 1'b0,x127 } )+$signed( -{ 1'b0,x383 } )+$signed( -{ 1'b0,x639 } )+$signed(11'd16);
assign y159=temp_y[159][11] ==1'b1 ? 5'd0 :  
        temp_y[159][8] ==1'b1 ? 5'd31 : 
        temp_y[159][2]==1'b1 ? temp_y[159][7:3]+1'b1 : temp_y[159][7:3];
assign temp_y[223] = 
+$signed( { 1'b0,x110 }  )+$signed( -{ 1'b0,x366 } )+$signed( { 1'b0,x111 }  )+$signed( -{ 1'b0,x367 } )+$signed( { 2'b0,x126 } <<<3'd1 )+$signed( -{ 1'b0,x382 } )+$signed( -{ 1'b0,x638 } )+$signed( { 2'b0,x127 } <<<3'd1 )+$signed( -{ 1'b0,x383 } )+$signed( -{ 2'b0,x639 }<<<3'd1 )+$signed(11'd40);
assign y223=temp_y[223][11] ==1'b1 ? 5'd0 :  
        temp_y[223][8] ==1'b1 ? 5'd31 : 
        temp_y[223][2]==1'b1 ? temp_y[223][7:3]+1'b1 : temp_y[223][7:3];
assign temp_y[287] = 
+$signed( -{ 1'b0,x110 } )+$signed( { 2'b0,x366 } <<<3'd1 )+$signed( -{ 1'b0,x622 } )+$signed( -{ 1'b0,x111 } )+$signed( { 2'b0,x367 } <<<3'd1 )+$signed( -{ 2'b0,x623 }<<<3'd1 )+$signed( -{ 1'b0,x126 } )+$signed( { 2'b0,x382 } <<<3'd1 )+$signed( -{ 1'b0,x638 } )+$signed( -{ 2'b0,x127 }<<<3'd1 )+$signed( { 3'b0,x383 }<<<3'd2 )+$signed( -{ 2'b0,x639 }<<<3'd1 )+$signed(11'd32);
assign y287=temp_y[287][11] ==1'b1 ? 5'd0 :  
        temp_y[287][8] ==1'b1 ? 5'd31 : 
        temp_y[287][2]==1'b1 ? temp_y[287][7:3]+1'b1 : temp_y[287][7:3];
assign temp_y[351] = 
+$signed( -{ 1'b0,x110 } )+$signed( -{ 2'b0,x366 }<<<3'd1 )+$signed( -{ 1'b0,x622 } )+$signed( { 1'b0,x111 }  )+$signed( { 2'b0,x367 } <<<3'd1 )+$signed( { 1'b0,x623 }  )+$signed( { 1'b0,x126 }  )+$signed( { 2'b0,x382 } <<<3'd1 )+$signed( { 2'b0,x638 } <<<3'd1 )+$signed( -{ 1'b0,x127 } )+$signed( -{ 2'b0,x383 }<<<3'd1 )+$signed( -{ 1'b0,x639 } )-$signed(11'd68);
assign y351=temp_y[351][11] ==1'b1 ? 5'd0 :  
        temp_y[351][8] ==1'b1 ? 5'd31 : 
        temp_y[351][2]==1'b1 ? temp_y[351][7:3]+1'b1 : temp_y[351][7:3];
assign temp_y[415] = 
+$signed( { 1'b0,x366 }  )+$signed( { 1'b0,x623 }  )+$signed( { 1'b0,x639 }  )-$signed(11'd108);
assign y415=temp_y[415][11] ==1'b1 ? 5'd0 :  
        temp_y[415][8] ==1'b1 ? 5'd31 : 
        temp_y[415][2]==1'b1 ? temp_y[415][7:3]+1'b1 : temp_y[415][7:3];
assign temp_y[479] = 
+$signed( -{ 2'b0,x110 }<<<3'd1 )+$signed( { 2'b0,x622 } <<<3'd1 )+$signed( -{ 2'b0,x111 }<<<3'd1 )+$signed( { 1'b0,x367 }  )+$signed( { 1'b0,x623 }  )+$signed( -{ 2'b0,x126 }<<<3'd1 )+$signed( { 1'b0,x382 }  )+$signed( { 1'b0,x638 }  )+$signed( -{ 1'b0,x127 } )+$signed(11'd64);
assign y479=temp_y[479][11] ==1'b1 ? 5'd0 :  
        temp_y[479][8] ==1'b1 ? 5'd31 : 
        temp_y[479][2]==1'b1 ? temp_y[479][7:3]+1'b1 : temp_y[479][7:3];
assign temp_y[543] = 
+$signed( -{ 2'b0,x110 }<<<3'd1 )+$signed( -{ 1'b0,x366 } )+$signed( -{ 3'b0,x111 }<<<3'd2)+$signed( { 1'b0,x126 }  )+$signed( { 1'b0,x382 }  )+$signed( { 3'b0,x127 }<<<3'd2 )+$signed(11'd16);
assign y543=temp_y[543][11] ==1'b1 ? 5'd0 :  
        temp_y[543][8] ==1'b1 ? 5'd31 : 
        temp_y[543][2]==1'b1 ? temp_y[543][7:3]+1'b1 : temp_y[543][7:3];
assign temp_y[607] = 
+$signed( { 2'b0,x366 } <<<3'd1 )+$signed( { 2'b0,x622 } <<<3'd1 )+$signed( -{ 1'b0,x111 } )+$signed( -{ 2'b0,x367 }<<<3'd1 )+$signed( -{ 2'b0,x623 }<<<3'd1 )+$signed( { 2'b0,x382 } <<<3'd1 )+$signed( { 1'b0,x638 }  )+$signed( -{ 2'b0,x383 }<<<3'd1 )-$signed(11'd8);
assign y607=temp_y[607][11] ==1'b1 ? 5'd0 :  
        temp_y[607][8] ==1'b1 ? 5'd31 : 
        temp_y[607][2]==1'b1 ? temp_y[607][7:3]+1'b1 : temp_y[607][7:3];
assign temp_y[32] = 
+$signed( -{ 2'b0,x384 }<<<3'd1 )+$signed( -{ 1'b0,x640 } )+$signed( { 1'b0,x129 }  )+$signed( { 1'b0,x385 }  )+$signed( { 1'b0,x641 }  )+$signed( -{ 2'b0,x400 }<<<3'd1 )+$signed( -{ 2'b0,x656 }<<<3'd1 )+$signed( { 2'b0,x401 } <<<3'd1 )+$signed( { 2'b0,x657 } <<<3'd1 )-$signed(11'd16);
assign y32=temp_y[32][11] ==1'b1 ? 5'd0 :  
        temp_y[32][8] ==1'b1 ? 5'd31 : 
        temp_y[32][2]==1'b1 ? temp_y[32][7:3]+1'b1 : temp_y[32][7:3];
assign temp_y[96] = 
+$signed( { 3'b0,x128 }<<<3'd2 )+$signed( -{ 2'b0,x384 }<<<3'd1 )+$signed( -{ 2'b0,x640 }<<<3'd1 )+$signed( { 2'b0,x129 } <<<3'd1 )+$signed( -{ 3'b0,x385 }<<<3'd2)+$signed( { 1'b0,x641 }  )+$signed( -{ 1'b0,x144 } )+$signed( { 1'b0,x656 }  )+$signed( -{ 2'b0,x145 }<<<3'd1 )+$signed( -{ 1'b0,x401 } )+$signed( { 2'b0,x657 } <<<3'd1 )+$signed(11'd24);
assign y96=temp_y[96][11] ==1'b1 ? 5'd0 :  
        temp_y[96][8] ==1'b1 ? 5'd31 : 
        temp_y[96][2]==1'b1 ? temp_y[96][7:3]+1'b1 : temp_y[96][7:3];
assign temp_y[160] = 
+$signed( { 2'b0,x128 } <<<3'd1 )+$signed( { 2'b0,x384 } <<<3'd1 )+$signed( { 1'b0,x640 }  )+$signed( { 2'b0,x129 } <<<3'd1 )+$signed( -{ 1'b0,x385 } )+$signed( { 1'b0,x641 }  )+$signed( -{ 2'b0,x144 }<<<3'd1 )+$signed( -{ 2'b0,x400 }<<<3'd1 )+$signed( -{ 1'b0,x656 } )+$signed( -{ 1'b0,x145 } )+$signed( -{ 1'b0,x401 } )+$signed( -{ 1'b0,x657 } )+$signed(11'd16);
assign y160=temp_y[160][11] ==1'b1 ? 5'd0 :  
        temp_y[160][8] ==1'b1 ? 5'd31 : 
        temp_y[160][2]==1'b1 ? temp_y[160][7:3]+1'b1 : temp_y[160][7:3];
assign temp_y[224] = 
+$signed( { 1'b0,x128 }  )+$signed( -{ 1'b0,x384 } )+$signed( { 1'b0,x129 }  )+$signed( -{ 1'b0,x385 } )+$signed( { 2'b0,x144 } <<<3'd1 )+$signed( -{ 1'b0,x400 } )+$signed( -{ 1'b0,x656 } )+$signed( { 2'b0,x145 } <<<3'd1 )+$signed( -{ 1'b0,x401 } )+$signed( -{ 2'b0,x657 }<<<3'd1 )+$signed(11'd40);
assign y224=temp_y[224][11] ==1'b1 ? 5'd0 :  
        temp_y[224][8] ==1'b1 ? 5'd31 : 
        temp_y[224][2]==1'b1 ? temp_y[224][7:3]+1'b1 : temp_y[224][7:3];
assign temp_y[288] = 
+$signed( -{ 1'b0,x128 } )+$signed( { 2'b0,x384 } <<<3'd1 )+$signed( -{ 1'b0,x640 } )+$signed( -{ 1'b0,x129 } )+$signed( { 2'b0,x385 } <<<3'd1 )+$signed( -{ 2'b0,x641 }<<<3'd1 )+$signed( -{ 1'b0,x144 } )+$signed( { 2'b0,x400 } <<<3'd1 )+$signed( -{ 1'b0,x656 } )+$signed( -{ 2'b0,x145 }<<<3'd1 )+$signed( { 3'b0,x401 }<<<3'd2 )+$signed( -{ 2'b0,x657 }<<<3'd1 )+$signed(11'd32);
assign y288=temp_y[288][11] ==1'b1 ? 5'd0 :  
        temp_y[288][8] ==1'b1 ? 5'd31 : 
        temp_y[288][2]==1'b1 ? temp_y[288][7:3]+1'b1 : temp_y[288][7:3];
assign temp_y[352] = 
+$signed( -{ 1'b0,x128 } )+$signed( -{ 2'b0,x384 }<<<3'd1 )+$signed( -{ 1'b0,x640 } )+$signed( { 1'b0,x129 }  )+$signed( { 2'b0,x385 } <<<3'd1 )+$signed( { 1'b0,x641 }  )+$signed( { 1'b0,x144 }  )+$signed( { 2'b0,x400 } <<<3'd1 )+$signed( { 2'b0,x656 } <<<3'd1 )+$signed( -{ 1'b0,x145 } )+$signed( -{ 2'b0,x401 }<<<3'd1 )+$signed( -{ 1'b0,x657 } )-$signed(11'd68);
assign y352=temp_y[352][11] ==1'b1 ? 5'd0 :  
        temp_y[352][8] ==1'b1 ? 5'd31 : 
        temp_y[352][2]==1'b1 ? temp_y[352][7:3]+1'b1 : temp_y[352][7:3];
assign temp_y[416] = 
+$signed( { 1'b0,x384 }  )+$signed( { 1'b0,x641 }  )+$signed( { 1'b0,x657 }  )-$signed(11'd108);
assign y416=temp_y[416][11] ==1'b1 ? 5'd0 :  
        temp_y[416][8] ==1'b1 ? 5'd31 : 
        temp_y[416][2]==1'b1 ? temp_y[416][7:3]+1'b1 : temp_y[416][7:3];
assign temp_y[480] = 
+$signed( -{ 2'b0,x128 }<<<3'd1 )+$signed( { 2'b0,x640 } <<<3'd1 )+$signed( -{ 2'b0,x129 }<<<3'd1 )+$signed( { 1'b0,x385 }  )+$signed( { 1'b0,x641 }  )+$signed( -{ 2'b0,x144 }<<<3'd1 )+$signed( { 1'b0,x400 }  )+$signed( { 1'b0,x656 }  )+$signed( -{ 1'b0,x145 } )+$signed(11'd64);
assign y480=temp_y[480][11] ==1'b1 ? 5'd0 :  
        temp_y[480][8] ==1'b1 ? 5'd31 : 
        temp_y[480][2]==1'b1 ? temp_y[480][7:3]+1'b1 : temp_y[480][7:3];
assign temp_y[544] = 
+$signed( -{ 2'b0,x128 }<<<3'd1 )+$signed( -{ 1'b0,x384 } )+$signed( -{ 3'b0,x129 }<<<3'd2)+$signed( { 1'b0,x144 }  )+$signed( { 1'b0,x400 }  )+$signed( { 3'b0,x145 }<<<3'd2 )+$signed(11'd16);
assign y544=temp_y[544][11] ==1'b1 ? 5'd0 :  
        temp_y[544][8] ==1'b1 ? 5'd31 : 
        temp_y[544][2]==1'b1 ? temp_y[544][7:3]+1'b1 : temp_y[544][7:3];
assign temp_y[608] = 
+$signed( { 2'b0,x384 } <<<3'd1 )+$signed( { 2'b0,x640 } <<<3'd1 )+$signed( -{ 1'b0,x129 } )+$signed( -{ 2'b0,x385 }<<<3'd1 )+$signed( -{ 2'b0,x641 }<<<3'd1 )+$signed( { 2'b0,x400 } <<<3'd1 )+$signed( { 1'b0,x656 }  )+$signed( -{ 2'b0,x401 }<<<3'd1 )-$signed(11'd8);
assign y608=temp_y[608][11] ==1'b1 ? 5'd0 :  
        temp_y[608][8] ==1'b1 ? 5'd31 : 
        temp_y[608][2]==1'b1 ? temp_y[608][7:3]+1'b1 : temp_y[608][7:3];
assign temp_y[33] = 
+$signed( -{ 2'b0,x386 }<<<3'd1 )+$signed( -{ 1'b0,x642 } )+$signed( { 1'b0,x131 }  )+$signed( { 1'b0,x387 }  )+$signed( { 1'b0,x643 }  )+$signed( -{ 2'b0,x402 }<<<3'd1 )+$signed( -{ 2'b0,x658 }<<<3'd1 )+$signed( { 2'b0,x403 } <<<3'd1 )+$signed( { 2'b0,x659 } <<<3'd1 )-$signed(11'd16);
assign y33=temp_y[33][11] ==1'b1 ? 5'd0 :  
        temp_y[33][8] ==1'b1 ? 5'd31 : 
        temp_y[33][2]==1'b1 ? temp_y[33][7:3]+1'b1 : temp_y[33][7:3];
assign temp_y[97] = 
+$signed( { 3'b0,x130 }<<<3'd2 )+$signed( -{ 2'b0,x386 }<<<3'd1 )+$signed( -{ 2'b0,x642 }<<<3'd1 )+$signed( { 2'b0,x131 } <<<3'd1 )+$signed( -{ 3'b0,x387 }<<<3'd2)+$signed( { 1'b0,x643 }  )+$signed( -{ 1'b0,x146 } )+$signed( { 1'b0,x658 }  )+$signed( -{ 2'b0,x147 }<<<3'd1 )+$signed( -{ 1'b0,x403 } )+$signed( { 2'b0,x659 } <<<3'd1 )+$signed(11'd24);
assign y97=temp_y[97][11] ==1'b1 ? 5'd0 :  
        temp_y[97][8] ==1'b1 ? 5'd31 : 
        temp_y[97][2]==1'b1 ? temp_y[97][7:3]+1'b1 : temp_y[97][7:3];
assign temp_y[161] = 
+$signed( { 2'b0,x130 } <<<3'd1 )+$signed( { 2'b0,x386 } <<<3'd1 )+$signed( { 1'b0,x642 }  )+$signed( { 2'b0,x131 } <<<3'd1 )+$signed( -{ 1'b0,x387 } )+$signed( { 1'b0,x643 }  )+$signed( -{ 2'b0,x146 }<<<3'd1 )+$signed( -{ 2'b0,x402 }<<<3'd1 )+$signed( -{ 1'b0,x658 } )+$signed( -{ 1'b0,x147 } )+$signed( -{ 1'b0,x403 } )+$signed( -{ 1'b0,x659 } )+$signed(11'd16);
assign y161=temp_y[161][11] ==1'b1 ? 5'd0 :  
        temp_y[161][8] ==1'b1 ? 5'd31 : 
        temp_y[161][2]==1'b1 ? temp_y[161][7:3]+1'b1 : temp_y[161][7:3];
assign temp_y[225] = 
+$signed( { 1'b0,x130 }  )+$signed( -{ 1'b0,x386 } )+$signed( { 1'b0,x131 }  )+$signed( -{ 1'b0,x387 } )+$signed( { 2'b0,x146 } <<<3'd1 )+$signed( -{ 1'b0,x402 } )+$signed( -{ 1'b0,x658 } )+$signed( { 2'b0,x147 } <<<3'd1 )+$signed( -{ 1'b0,x403 } )+$signed( -{ 2'b0,x659 }<<<3'd1 )+$signed(11'd40);
assign y225=temp_y[225][11] ==1'b1 ? 5'd0 :  
        temp_y[225][8] ==1'b1 ? 5'd31 : 
        temp_y[225][2]==1'b1 ? temp_y[225][7:3]+1'b1 : temp_y[225][7:3];
assign temp_y[289] = 
+$signed( -{ 1'b0,x130 } )+$signed( { 2'b0,x386 } <<<3'd1 )+$signed( -{ 1'b0,x642 } )+$signed( -{ 1'b0,x131 } )+$signed( { 2'b0,x387 } <<<3'd1 )+$signed( -{ 2'b0,x643 }<<<3'd1 )+$signed( -{ 1'b0,x146 } )+$signed( { 2'b0,x402 } <<<3'd1 )+$signed( -{ 1'b0,x658 } )+$signed( -{ 2'b0,x147 }<<<3'd1 )+$signed( { 3'b0,x403 }<<<3'd2 )+$signed( -{ 2'b0,x659 }<<<3'd1 )+$signed(11'd32);
assign y289=temp_y[289][11] ==1'b1 ? 5'd0 :  
        temp_y[289][8] ==1'b1 ? 5'd31 : 
        temp_y[289][2]==1'b1 ? temp_y[289][7:3]+1'b1 : temp_y[289][7:3];
assign temp_y[353] = 
+$signed( -{ 1'b0,x130 } )+$signed( -{ 2'b0,x386 }<<<3'd1 )+$signed( -{ 1'b0,x642 } )+$signed( { 1'b0,x131 }  )+$signed( { 2'b0,x387 } <<<3'd1 )+$signed( { 1'b0,x643 }  )+$signed( { 1'b0,x146 }  )+$signed( { 2'b0,x402 } <<<3'd1 )+$signed( { 2'b0,x658 } <<<3'd1 )+$signed( -{ 1'b0,x147 } )+$signed( -{ 2'b0,x403 }<<<3'd1 )+$signed( -{ 1'b0,x659 } )-$signed(11'd68);
assign y353=temp_y[353][11] ==1'b1 ? 5'd0 :  
        temp_y[353][8] ==1'b1 ? 5'd31 : 
        temp_y[353][2]==1'b1 ? temp_y[353][7:3]+1'b1 : temp_y[353][7:3];
assign temp_y[417] = 
+$signed( { 1'b0,x386 }  )+$signed( { 1'b0,x643 }  )+$signed( { 1'b0,x659 }  )-$signed(11'd108);
assign y417=temp_y[417][11] ==1'b1 ? 5'd0 :  
        temp_y[417][8] ==1'b1 ? 5'd31 : 
        temp_y[417][2]==1'b1 ? temp_y[417][7:3]+1'b1 : temp_y[417][7:3];
assign temp_y[481] = 
+$signed( -{ 2'b0,x130 }<<<3'd1 )+$signed( { 2'b0,x642 } <<<3'd1 )+$signed( -{ 2'b0,x131 }<<<3'd1 )+$signed( { 1'b0,x387 }  )+$signed( { 1'b0,x643 }  )+$signed( -{ 2'b0,x146 }<<<3'd1 )+$signed( { 1'b0,x402 }  )+$signed( { 1'b0,x658 }  )+$signed( -{ 1'b0,x147 } )+$signed(11'd64);
assign y481=temp_y[481][11] ==1'b1 ? 5'd0 :  
        temp_y[481][8] ==1'b1 ? 5'd31 : 
        temp_y[481][2]==1'b1 ? temp_y[481][7:3]+1'b1 : temp_y[481][7:3];
assign temp_y[545] = 
+$signed( -{ 2'b0,x130 }<<<3'd1 )+$signed( -{ 1'b0,x386 } )+$signed( -{ 3'b0,x131 }<<<3'd2)+$signed( { 1'b0,x146 }  )+$signed( { 1'b0,x402 }  )+$signed( { 3'b0,x147 }<<<3'd2 )+$signed(11'd16);
assign y545=temp_y[545][11] ==1'b1 ? 5'd0 :  
        temp_y[545][8] ==1'b1 ? 5'd31 : 
        temp_y[545][2]==1'b1 ? temp_y[545][7:3]+1'b1 : temp_y[545][7:3];
assign temp_y[609] = 
+$signed( { 2'b0,x386 } <<<3'd1 )+$signed( { 2'b0,x642 } <<<3'd1 )+$signed( -{ 1'b0,x131 } )+$signed( -{ 2'b0,x387 }<<<3'd1 )+$signed( -{ 2'b0,x643 }<<<3'd1 )+$signed( { 2'b0,x402 } <<<3'd1 )+$signed( { 1'b0,x658 }  )+$signed( -{ 2'b0,x403 }<<<3'd1 )-$signed(11'd8);
assign y609=temp_y[609][11] ==1'b1 ? 5'd0 :  
        temp_y[609][8] ==1'b1 ? 5'd31 : 
        temp_y[609][2]==1'b1 ? temp_y[609][7:3]+1'b1 : temp_y[609][7:3];
assign temp_y[34] = 
+$signed( -{ 2'b0,x388 }<<<3'd1 )+$signed( -{ 1'b0,x644 } )+$signed( { 1'b0,x133 }  )+$signed( { 1'b0,x389 }  )+$signed( { 1'b0,x645 }  )+$signed( -{ 2'b0,x404 }<<<3'd1 )+$signed( -{ 2'b0,x660 }<<<3'd1 )+$signed( { 2'b0,x405 } <<<3'd1 )+$signed( { 2'b0,x661 } <<<3'd1 )-$signed(11'd16);
assign y34=temp_y[34][11] ==1'b1 ? 5'd0 :  
        temp_y[34][8] ==1'b1 ? 5'd31 : 
        temp_y[34][2]==1'b1 ? temp_y[34][7:3]+1'b1 : temp_y[34][7:3];
assign temp_y[98] = 
+$signed( { 3'b0,x132 }<<<3'd2 )+$signed( -{ 2'b0,x388 }<<<3'd1 )+$signed( -{ 2'b0,x644 }<<<3'd1 )+$signed( { 2'b0,x133 } <<<3'd1 )+$signed( -{ 3'b0,x389 }<<<3'd2)+$signed( { 1'b0,x645 }  )+$signed( -{ 1'b0,x148 } )+$signed( { 1'b0,x660 }  )+$signed( -{ 2'b0,x149 }<<<3'd1 )+$signed( -{ 1'b0,x405 } )+$signed( { 2'b0,x661 } <<<3'd1 )+$signed(11'd24);
assign y98=temp_y[98][11] ==1'b1 ? 5'd0 :  
        temp_y[98][8] ==1'b1 ? 5'd31 : 
        temp_y[98][2]==1'b1 ? temp_y[98][7:3]+1'b1 : temp_y[98][7:3];
assign temp_y[162] = 
+$signed( { 2'b0,x132 } <<<3'd1 )+$signed( { 2'b0,x388 } <<<3'd1 )+$signed( { 1'b0,x644 }  )+$signed( { 2'b0,x133 } <<<3'd1 )+$signed( -{ 1'b0,x389 } )+$signed( { 1'b0,x645 }  )+$signed( -{ 2'b0,x148 }<<<3'd1 )+$signed( -{ 2'b0,x404 }<<<3'd1 )+$signed( -{ 1'b0,x660 } )+$signed( -{ 1'b0,x149 } )+$signed( -{ 1'b0,x405 } )+$signed( -{ 1'b0,x661 } )+$signed(11'd16);
assign y162=temp_y[162][11] ==1'b1 ? 5'd0 :  
        temp_y[162][8] ==1'b1 ? 5'd31 : 
        temp_y[162][2]==1'b1 ? temp_y[162][7:3]+1'b1 : temp_y[162][7:3];
assign temp_y[226] = 
+$signed( { 1'b0,x132 }  )+$signed( -{ 1'b0,x388 } )+$signed( { 1'b0,x133 }  )+$signed( -{ 1'b0,x389 } )+$signed( { 2'b0,x148 } <<<3'd1 )+$signed( -{ 1'b0,x404 } )+$signed( -{ 1'b0,x660 } )+$signed( { 2'b0,x149 } <<<3'd1 )+$signed( -{ 1'b0,x405 } )+$signed( -{ 2'b0,x661 }<<<3'd1 )+$signed(11'd40);
assign y226=temp_y[226][11] ==1'b1 ? 5'd0 :  
        temp_y[226][8] ==1'b1 ? 5'd31 : 
        temp_y[226][2]==1'b1 ? temp_y[226][7:3]+1'b1 : temp_y[226][7:3];
assign temp_y[290] = 
+$signed( -{ 1'b0,x132 } )+$signed( { 2'b0,x388 } <<<3'd1 )+$signed( -{ 1'b0,x644 } )+$signed( -{ 1'b0,x133 } )+$signed( { 2'b0,x389 } <<<3'd1 )+$signed( -{ 2'b0,x645 }<<<3'd1 )+$signed( -{ 1'b0,x148 } )+$signed( { 2'b0,x404 } <<<3'd1 )+$signed( -{ 1'b0,x660 } )+$signed( -{ 2'b0,x149 }<<<3'd1 )+$signed( { 3'b0,x405 }<<<3'd2 )+$signed( -{ 2'b0,x661 }<<<3'd1 )+$signed(11'd32);
assign y290=temp_y[290][11] ==1'b1 ? 5'd0 :  
        temp_y[290][8] ==1'b1 ? 5'd31 : 
        temp_y[290][2]==1'b1 ? temp_y[290][7:3]+1'b1 : temp_y[290][7:3];
assign temp_y[354] = 
+$signed( -{ 1'b0,x132 } )+$signed( -{ 2'b0,x388 }<<<3'd1 )+$signed( -{ 1'b0,x644 } )+$signed( { 1'b0,x133 }  )+$signed( { 2'b0,x389 } <<<3'd1 )+$signed( { 1'b0,x645 }  )+$signed( { 1'b0,x148 }  )+$signed( { 2'b0,x404 } <<<3'd1 )+$signed( { 2'b0,x660 } <<<3'd1 )+$signed( -{ 1'b0,x149 } )+$signed( -{ 2'b0,x405 }<<<3'd1 )+$signed( -{ 1'b0,x661 } )-$signed(11'd68);
assign y354=temp_y[354][11] ==1'b1 ? 5'd0 :  
        temp_y[354][8] ==1'b1 ? 5'd31 : 
        temp_y[354][2]==1'b1 ? temp_y[354][7:3]+1'b1 : temp_y[354][7:3];
assign temp_y[418] = 
+$signed( { 1'b0,x388 }  )+$signed( { 1'b0,x645 }  )+$signed( { 1'b0,x661 }  )-$signed(11'd108);
assign y418=temp_y[418][11] ==1'b1 ? 5'd0 :  
        temp_y[418][8] ==1'b1 ? 5'd31 : 
        temp_y[418][2]==1'b1 ? temp_y[418][7:3]+1'b1 : temp_y[418][7:3];
assign temp_y[482] = 
+$signed( -{ 2'b0,x132 }<<<3'd1 )+$signed( { 2'b0,x644 } <<<3'd1 )+$signed( -{ 2'b0,x133 }<<<3'd1 )+$signed( { 1'b0,x389 }  )+$signed( { 1'b0,x645 }  )+$signed( -{ 2'b0,x148 }<<<3'd1 )+$signed( { 1'b0,x404 }  )+$signed( { 1'b0,x660 }  )+$signed( -{ 1'b0,x149 } )+$signed(11'd64);
assign y482=temp_y[482][11] ==1'b1 ? 5'd0 :  
        temp_y[482][8] ==1'b1 ? 5'd31 : 
        temp_y[482][2]==1'b1 ? temp_y[482][7:3]+1'b1 : temp_y[482][7:3];
assign temp_y[546] = 
+$signed( -{ 2'b0,x132 }<<<3'd1 )+$signed( -{ 1'b0,x388 } )+$signed( -{ 3'b0,x133 }<<<3'd2)+$signed( { 1'b0,x148 }  )+$signed( { 1'b0,x404 }  )+$signed( { 3'b0,x149 }<<<3'd2 )+$signed(11'd16);
assign y546=temp_y[546][11] ==1'b1 ? 5'd0 :  
        temp_y[546][8] ==1'b1 ? 5'd31 : 
        temp_y[546][2]==1'b1 ? temp_y[546][7:3]+1'b1 : temp_y[546][7:3];
assign temp_y[610] = 
+$signed( { 2'b0,x388 } <<<3'd1 )+$signed( { 2'b0,x644 } <<<3'd1 )+$signed( -{ 1'b0,x133 } )+$signed( -{ 2'b0,x389 }<<<3'd1 )+$signed( -{ 2'b0,x645 }<<<3'd1 )+$signed( { 2'b0,x404 } <<<3'd1 )+$signed( { 1'b0,x660 }  )+$signed( -{ 2'b0,x405 }<<<3'd1 )-$signed(11'd8);
assign y610=temp_y[610][11] ==1'b1 ? 5'd0 :  
        temp_y[610][8] ==1'b1 ? 5'd31 : 
        temp_y[610][2]==1'b1 ? temp_y[610][7:3]+1'b1 : temp_y[610][7:3];
assign temp_y[35] = 
+$signed( -{ 2'b0,x390 }<<<3'd1 )+$signed( -{ 1'b0,x646 } )+$signed( { 1'b0,x135 }  )+$signed( { 1'b0,x391 }  )+$signed( { 1'b0,x647 }  )+$signed( -{ 2'b0,x406 }<<<3'd1 )+$signed( -{ 2'b0,x662 }<<<3'd1 )+$signed( { 2'b0,x407 } <<<3'd1 )+$signed( { 2'b0,x663 } <<<3'd1 )-$signed(11'd16);
assign y35=temp_y[35][11] ==1'b1 ? 5'd0 :  
        temp_y[35][8] ==1'b1 ? 5'd31 : 
        temp_y[35][2]==1'b1 ? temp_y[35][7:3]+1'b1 : temp_y[35][7:3];
assign temp_y[99] = 
+$signed( { 3'b0,x134 }<<<3'd2 )+$signed( -{ 2'b0,x390 }<<<3'd1 )+$signed( -{ 2'b0,x646 }<<<3'd1 )+$signed( { 2'b0,x135 } <<<3'd1 )+$signed( -{ 3'b0,x391 }<<<3'd2)+$signed( { 1'b0,x647 }  )+$signed( -{ 1'b0,x150 } )+$signed( { 1'b0,x662 }  )+$signed( -{ 2'b0,x151 }<<<3'd1 )+$signed( -{ 1'b0,x407 } )+$signed( { 2'b0,x663 } <<<3'd1 )+$signed(11'd24);
assign y99=temp_y[99][11] ==1'b1 ? 5'd0 :  
        temp_y[99][8] ==1'b1 ? 5'd31 : 
        temp_y[99][2]==1'b1 ? temp_y[99][7:3]+1'b1 : temp_y[99][7:3];
assign temp_y[163] = 
+$signed( { 2'b0,x134 } <<<3'd1 )+$signed( { 2'b0,x390 } <<<3'd1 )+$signed( { 1'b0,x646 }  )+$signed( { 2'b0,x135 } <<<3'd1 )+$signed( -{ 1'b0,x391 } )+$signed( { 1'b0,x647 }  )+$signed( -{ 2'b0,x150 }<<<3'd1 )+$signed( -{ 2'b0,x406 }<<<3'd1 )+$signed( -{ 1'b0,x662 } )+$signed( -{ 1'b0,x151 } )+$signed( -{ 1'b0,x407 } )+$signed( -{ 1'b0,x663 } )+$signed(11'd16);
assign y163=temp_y[163][11] ==1'b1 ? 5'd0 :  
        temp_y[163][8] ==1'b1 ? 5'd31 : 
        temp_y[163][2]==1'b1 ? temp_y[163][7:3]+1'b1 : temp_y[163][7:3];
assign temp_y[227] = 
+$signed( { 1'b0,x134 }  )+$signed( -{ 1'b0,x390 } )+$signed( { 1'b0,x135 }  )+$signed( -{ 1'b0,x391 } )+$signed( { 2'b0,x150 } <<<3'd1 )+$signed( -{ 1'b0,x406 } )+$signed( -{ 1'b0,x662 } )+$signed( { 2'b0,x151 } <<<3'd1 )+$signed( -{ 1'b0,x407 } )+$signed( -{ 2'b0,x663 }<<<3'd1 )+$signed(11'd40);
assign y227=temp_y[227][11] ==1'b1 ? 5'd0 :  
        temp_y[227][8] ==1'b1 ? 5'd31 : 
        temp_y[227][2]==1'b1 ? temp_y[227][7:3]+1'b1 : temp_y[227][7:3];
assign temp_y[291] = 
+$signed( -{ 1'b0,x134 } )+$signed( { 2'b0,x390 } <<<3'd1 )+$signed( -{ 1'b0,x646 } )+$signed( -{ 1'b0,x135 } )+$signed( { 2'b0,x391 } <<<3'd1 )+$signed( -{ 2'b0,x647 }<<<3'd1 )+$signed( -{ 1'b0,x150 } )+$signed( { 2'b0,x406 } <<<3'd1 )+$signed( -{ 1'b0,x662 } )+$signed( -{ 2'b0,x151 }<<<3'd1 )+$signed( { 3'b0,x407 }<<<3'd2 )+$signed( -{ 2'b0,x663 }<<<3'd1 )+$signed(11'd32);
assign y291=temp_y[291][11] ==1'b1 ? 5'd0 :  
        temp_y[291][8] ==1'b1 ? 5'd31 : 
        temp_y[291][2]==1'b1 ? temp_y[291][7:3]+1'b1 : temp_y[291][7:3];
assign temp_y[355] = 
+$signed( -{ 1'b0,x134 } )+$signed( -{ 2'b0,x390 }<<<3'd1 )+$signed( -{ 1'b0,x646 } )+$signed( { 1'b0,x135 }  )+$signed( { 2'b0,x391 } <<<3'd1 )+$signed( { 1'b0,x647 }  )+$signed( { 1'b0,x150 }  )+$signed( { 2'b0,x406 } <<<3'd1 )+$signed( { 2'b0,x662 } <<<3'd1 )+$signed( -{ 1'b0,x151 } )+$signed( -{ 2'b0,x407 }<<<3'd1 )+$signed( -{ 1'b0,x663 } )-$signed(11'd68);
assign y355=temp_y[355][11] ==1'b1 ? 5'd0 :  
        temp_y[355][8] ==1'b1 ? 5'd31 : 
        temp_y[355][2]==1'b1 ? temp_y[355][7:3]+1'b1 : temp_y[355][7:3];
assign temp_y[419] = 
+$signed( { 1'b0,x390 }  )+$signed( { 1'b0,x647 }  )+$signed( { 1'b0,x663 }  )-$signed(11'd108);
assign y419=temp_y[419][11] ==1'b1 ? 5'd0 :  
        temp_y[419][8] ==1'b1 ? 5'd31 : 
        temp_y[419][2]==1'b1 ? temp_y[419][7:3]+1'b1 : temp_y[419][7:3];
assign temp_y[483] = 
+$signed( -{ 2'b0,x134 }<<<3'd1 )+$signed( { 2'b0,x646 } <<<3'd1 )+$signed( -{ 2'b0,x135 }<<<3'd1 )+$signed( { 1'b0,x391 }  )+$signed( { 1'b0,x647 }  )+$signed( -{ 2'b0,x150 }<<<3'd1 )+$signed( { 1'b0,x406 }  )+$signed( { 1'b0,x662 }  )+$signed( -{ 1'b0,x151 } )+$signed(11'd64);
assign y483=temp_y[483][11] ==1'b1 ? 5'd0 :  
        temp_y[483][8] ==1'b1 ? 5'd31 : 
        temp_y[483][2]==1'b1 ? temp_y[483][7:3]+1'b1 : temp_y[483][7:3];
assign temp_y[547] = 
+$signed( -{ 2'b0,x134 }<<<3'd1 )+$signed( -{ 1'b0,x390 } )+$signed( -{ 3'b0,x135 }<<<3'd2)+$signed( { 1'b0,x150 }  )+$signed( { 1'b0,x406 }  )+$signed( { 3'b0,x151 }<<<3'd2 )+$signed(11'd16);
assign y547=temp_y[547][11] ==1'b1 ? 5'd0 :  
        temp_y[547][8] ==1'b1 ? 5'd31 : 
        temp_y[547][2]==1'b1 ? temp_y[547][7:3]+1'b1 : temp_y[547][7:3];
assign temp_y[611] = 
+$signed( { 2'b0,x390 } <<<3'd1 )+$signed( { 2'b0,x646 } <<<3'd1 )+$signed( -{ 1'b0,x135 } )+$signed( -{ 2'b0,x391 }<<<3'd1 )+$signed( -{ 2'b0,x647 }<<<3'd1 )+$signed( { 2'b0,x406 } <<<3'd1 )+$signed( { 1'b0,x662 }  )+$signed( -{ 2'b0,x407 }<<<3'd1 )-$signed(11'd8);
assign y611=temp_y[611][11] ==1'b1 ? 5'd0 :  
        temp_y[611][8] ==1'b1 ? 5'd31 : 
        temp_y[611][2]==1'b1 ? temp_y[611][7:3]+1'b1 : temp_y[611][7:3];
assign temp_y[36] = 
+$signed( -{ 2'b0,x392 }<<<3'd1 )+$signed( -{ 1'b0,x648 } )+$signed( { 1'b0,x137 }  )+$signed( { 1'b0,x393 }  )+$signed( { 1'b0,x649 }  )+$signed( -{ 2'b0,x408 }<<<3'd1 )+$signed( -{ 2'b0,x664 }<<<3'd1 )+$signed( { 2'b0,x409 } <<<3'd1 )+$signed( { 2'b0,x665 } <<<3'd1 )-$signed(11'd16);
assign y36=temp_y[36][11] ==1'b1 ? 5'd0 :  
        temp_y[36][8] ==1'b1 ? 5'd31 : 
        temp_y[36][2]==1'b1 ? temp_y[36][7:3]+1'b1 : temp_y[36][7:3];
assign temp_y[100] = 
+$signed( { 3'b0,x136 }<<<3'd2 )+$signed( -{ 2'b0,x392 }<<<3'd1 )+$signed( -{ 2'b0,x648 }<<<3'd1 )+$signed( { 2'b0,x137 } <<<3'd1 )+$signed( -{ 3'b0,x393 }<<<3'd2)+$signed( { 1'b0,x649 }  )+$signed( -{ 1'b0,x152 } )+$signed( { 1'b0,x664 }  )+$signed( -{ 2'b0,x153 }<<<3'd1 )+$signed( -{ 1'b0,x409 } )+$signed( { 2'b0,x665 } <<<3'd1 )+$signed(11'd24);
assign y100=temp_y[100][11] ==1'b1 ? 5'd0 :  
        temp_y[100][8] ==1'b1 ? 5'd31 : 
        temp_y[100][2]==1'b1 ? temp_y[100][7:3]+1'b1 : temp_y[100][7:3];
assign temp_y[164] = 
+$signed( { 2'b0,x136 } <<<3'd1 )+$signed( { 2'b0,x392 } <<<3'd1 )+$signed( { 1'b0,x648 }  )+$signed( { 2'b0,x137 } <<<3'd1 )+$signed( -{ 1'b0,x393 } )+$signed( { 1'b0,x649 }  )+$signed( -{ 2'b0,x152 }<<<3'd1 )+$signed( -{ 2'b0,x408 }<<<3'd1 )+$signed( -{ 1'b0,x664 } )+$signed( -{ 1'b0,x153 } )+$signed( -{ 1'b0,x409 } )+$signed( -{ 1'b0,x665 } )+$signed(11'd16);
assign y164=temp_y[164][11] ==1'b1 ? 5'd0 :  
        temp_y[164][8] ==1'b1 ? 5'd31 : 
        temp_y[164][2]==1'b1 ? temp_y[164][7:3]+1'b1 : temp_y[164][7:3];
assign temp_y[228] = 
+$signed( { 1'b0,x136 }  )+$signed( -{ 1'b0,x392 } )+$signed( { 1'b0,x137 }  )+$signed( -{ 1'b0,x393 } )+$signed( { 2'b0,x152 } <<<3'd1 )+$signed( -{ 1'b0,x408 } )+$signed( -{ 1'b0,x664 } )+$signed( { 2'b0,x153 } <<<3'd1 )+$signed( -{ 1'b0,x409 } )+$signed( -{ 2'b0,x665 }<<<3'd1 )+$signed(11'd40);
assign y228=temp_y[228][11] ==1'b1 ? 5'd0 :  
        temp_y[228][8] ==1'b1 ? 5'd31 : 
        temp_y[228][2]==1'b1 ? temp_y[228][7:3]+1'b1 : temp_y[228][7:3];
assign temp_y[292] = 
+$signed( -{ 1'b0,x136 } )+$signed( { 2'b0,x392 } <<<3'd1 )+$signed( -{ 1'b0,x648 } )+$signed( -{ 1'b0,x137 } )+$signed( { 2'b0,x393 } <<<3'd1 )+$signed( -{ 2'b0,x649 }<<<3'd1 )+$signed( -{ 1'b0,x152 } )+$signed( { 2'b0,x408 } <<<3'd1 )+$signed( -{ 1'b0,x664 } )+$signed( -{ 2'b0,x153 }<<<3'd1 )+$signed( { 3'b0,x409 }<<<3'd2 )+$signed( -{ 2'b0,x665 }<<<3'd1 )+$signed(11'd32);
assign y292=temp_y[292][11] ==1'b1 ? 5'd0 :  
        temp_y[292][8] ==1'b1 ? 5'd31 : 
        temp_y[292][2]==1'b1 ? temp_y[292][7:3]+1'b1 : temp_y[292][7:3];
assign temp_y[356] = 
+$signed( -{ 1'b0,x136 } )+$signed( -{ 2'b0,x392 }<<<3'd1 )+$signed( -{ 1'b0,x648 } )+$signed( { 1'b0,x137 }  )+$signed( { 2'b0,x393 } <<<3'd1 )+$signed( { 1'b0,x649 }  )+$signed( { 1'b0,x152 }  )+$signed( { 2'b0,x408 } <<<3'd1 )+$signed( { 2'b0,x664 } <<<3'd1 )+$signed( -{ 1'b0,x153 } )+$signed( -{ 2'b0,x409 }<<<3'd1 )+$signed( -{ 1'b0,x665 } )-$signed(11'd68);
assign y356=temp_y[356][11] ==1'b1 ? 5'd0 :  
        temp_y[356][8] ==1'b1 ? 5'd31 : 
        temp_y[356][2]==1'b1 ? temp_y[356][7:3]+1'b1 : temp_y[356][7:3];
assign temp_y[420] = 
+$signed( { 1'b0,x392 }  )+$signed( { 1'b0,x649 }  )+$signed( { 1'b0,x665 }  )-$signed(11'd108);
assign y420=temp_y[420][11] ==1'b1 ? 5'd0 :  
        temp_y[420][8] ==1'b1 ? 5'd31 : 
        temp_y[420][2]==1'b1 ? temp_y[420][7:3]+1'b1 : temp_y[420][7:3];
assign temp_y[484] = 
+$signed( -{ 2'b0,x136 }<<<3'd1 )+$signed( { 2'b0,x648 } <<<3'd1 )+$signed( -{ 2'b0,x137 }<<<3'd1 )+$signed( { 1'b0,x393 }  )+$signed( { 1'b0,x649 }  )+$signed( -{ 2'b0,x152 }<<<3'd1 )+$signed( { 1'b0,x408 }  )+$signed( { 1'b0,x664 }  )+$signed( -{ 1'b0,x153 } )+$signed(11'd64);
assign y484=temp_y[484][11] ==1'b1 ? 5'd0 :  
        temp_y[484][8] ==1'b1 ? 5'd31 : 
        temp_y[484][2]==1'b1 ? temp_y[484][7:3]+1'b1 : temp_y[484][7:3];
assign temp_y[548] = 
+$signed( -{ 2'b0,x136 }<<<3'd1 )+$signed( -{ 1'b0,x392 } )+$signed( -{ 3'b0,x137 }<<<3'd2)+$signed( { 1'b0,x152 }  )+$signed( { 1'b0,x408 }  )+$signed( { 3'b0,x153 }<<<3'd2 )+$signed(11'd16);
assign y548=temp_y[548][11] ==1'b1 ? 5'd0 :  
        temp_y[548][8] ==1'b1 ? 5'd31 : 
        temp_y[548][2]==1'b1 ? temp_y[548][7:3]+1'b1 : temp_y[548][7:3];
assign temp_y[612] = 
+$signed( { 2'b0,x392 } <<<3'd1 )+$signed( { 2'b0,x648 } <<<3'd1 )+$signed( -{ 1'b0,x137 } )+$signed( -{ 2'b0,x393 }<<<3'd1 )+$signed( -{ 2'b0,x649 }<<<3'd1 )+$signed( { 2'b0,x408 } <<<3'd1 )+$signed( { 1'b0,x664 }  )+$signed( -{ 2'b0,x409 }<<<3'd1 )-$signed(11'd8);
assign y612=temp_y[612][11] ==1'b1 ? 5'd0 :  
        temp_y[612][8] ==1'b1 ? 5'd31 : 
        temp_y[612][2]==1'b1 ? temp_y[612][7:3]+1'b1 : temp_y[612][7:3];
assign temp_y[37] = 
+$signed( -{ 2'b0,x394 }<<<3'd1 )+$signed( -{ 1'b0,x650 } )+$signed( { 1'b0,x139 }  )+$signed( { 1'b0,x395 }  )+$signed( { 1'b0,x651 }  )+$signed( -{ 2'b0,x410 }<<<3'd1 )+$signed( -{ 2'b0,x666 }<<<3'd1 )+$signed( { 2'b0,x411 } <<<3'd1 )+$signed( { 2'b0,x667 } <<<3'd1 )-$signed(11'd16);
assign y37=temp_y[37][11] ==1'b1 ? 5'd0 :  
        temp_y[37][8] ==1'b1 ? 5'd31 : 
        temp_y[37][2]==1'b1 ? temp_y[37][7:3]+1'b1 : temp_y[37][7:3];
assign temp_y[101] = 
+$signed( { 3'b0,x138 }<<<3'd2 )+$signed( -{ 2'b0,x394 }<<<3'd1 )+$signed( -{ 2'b0,x650 }<<<3'd1 )+$signed( { 2'b0,x139 } <<<3'd1 )+$signed( -{ 3'b0,x395 }<<<3'd2)+$signed( { 1'b0,x651 }  )+$signed( -{ 1'b0,x154 } )+$signed( { 1'b0,x666 }  )+$signed( -{ 2'b0,x155 }<<<3'd1 )+$signed( -{ 1'b0,x411 } )+$signed( { 2'b0,x667 } <<<3'd1 )+$signed(11'd24);
assign y101=temp_y[101][11] ==1'b1 ? 5'd0 :  
        temp_y[101][8] ==1'b1 ? 5'd31 : 
        temp_y[101][2]==1'b1 ? temp_y[101][7:3]+1'b1 : temp_y[101][7:3];
assign temp_y[165] = 
+$signed( { 2'b0,x138 } <<<3'd1 )+$signed( { 2'b0,x394 } <<<3'd1 )+$signed( { 1'b0,x650 }  )+$signed( { 2'b0,x139 } <<<3'd1 )+$signed( -{ 1'b0,x395 } )+$signed( { 1'b0,x651 }  )+$signed( -{ 2'b0,x154 }<<<3'd1 )+$signed( -{ 2'b0,x410 }<<<3'd1 )+$signed( -{ 1'b0,x666 } )+$signed( -{ 1'b0,x155 } )+$signed( -{ 1'b0,x411 } )+$signed( -{ 1'b0,x667 } )+$signed(11'd16);
assign y165=temp_y[165][11] ==1'b1 ? 5'd0 :  
        temp_y[165][8] ==1'b1 ? 5'd31 : 
        temp_y[165][2]==1'b1 ? temp_y[165][7:3]+1'b1 : temp_y[165][7:3];
assign temp_y[229] = 
+$signed( { 1'b0,x138 }  )+$signed( -{ 1'b0,x394 } )+$signed( { 1'b0,x139 }  )+$signed( -{ 1'b0,x395 } )+$signed( { 2'b0,x154 } <<<3'd1 )+$signed( -{ 1'b0,x410 } )+$signed( -{ 1'b0,x666 } )+$signed( { 2'b0,x155 } <<<3'd1 )+$signed( -{ 1'b0,x411 } )+$signed( -{ 2'b0,x667 }<<<3'd1 )+$signed(11'd40);
assign y229=temp_y[229][11] ==1'b1 ? 5'd0 :  
        temp_y[229][8] ==1'b1 ? 5'd31 : 
        temp_y[229][2]==1'b1 ? temp_y[229][7:3]+1'b1 : temp_y[229][7:3];
assign temp_y[293] = 
+$signed( -{ 1'b0,x138 } )+$signed( { 2'b0,x394 } <<<3'd1 )+$signed( -{ 1'b0,x650 } )+$signed( -{ 1'b0,x139 } )+$signed( { 2'b0,x395 } <<<3'd1 )+$signed( -{ 2'b0,x651 }<<<3'd1 )+$signed( -{ 1'b0,x154 } )+$signed( { 2'b0,x410 } <<<3'd1 )+$signed( -{ 1'b0,x666 } )+$signed( -{ 2'b0,x155 }<<<3'd1 )+$signed( { 3'b0,x411 }<<<3'd2 )+$signed( -{ 2'b0,x667 }<<<3'd1 )+$signed(11'd32);
assign y293=temp_y[293][11] ==1'b1 ? 5'd0 :  
        temp_y[293][8] ==1'b1 ? 5'd31 : 
        temp_y[293][2]==1'b1 ? temp_y[293][7:3]+1'b1 : temp_y[293][7:3];
assign temp_y[357] = 
+$signed( -{ 1'b0,x138 } )+$signed( -{ 2'b0,x394 }<<<3'd1 )+$signed( -{ 1'b0,x650 } )+$signed( { 1'b0,x139 }  )+$signed( { 2'b0,x395 } <<<3'd1 )+$signed( { 1'b0,x651 }  )+$signed( { 1'b0,x154 }  )+$signed( { 2'b0,x410 } <<<3'd1 )+$signed( { 2'b0,x666 } <<<3'd1 )+$signed( -{ 1'b0,x155 } )+$signed( -{ 2'b0,x411 }<<<3'd1 )+$signed( -{ 1'b0,x667 } )-$signed(11'd68);
assign y357=temp_y[357][11] ==1'b1 ? 5'd0 :  
        temp_y[357][8] ==1'b1 ? 5'd31 : 
        temp_y[357][2]==1'b1 ? temp_y[357][7:3]+1'b1 : temp_y[357][7:3];
assign temp_y[421] = 
+$signed( { 1'b0,x394 }  )+$signed( { 1'b0,x651 }  )+$signed( { 1'b0,x667 }  )-$signed(11'd108);
assign y421=temp_y[421][11] ==1'b1 ? 5'd0 :  
        temp_y[421][8] ==1'b1 ? 5'd31 : 
        temp_y[421][2]==1'b1 ? temp_y[421][7:3]+1'b1 : temp_y[421][7:3];
assign temp_y[485] = 
+$signed( -{ 2'b0,x138 }<<<3'd1 )+$signed( { 2'b0,x650 } <<<3'd1 )+$signed( -{ 2'b0,x139 }<<<3'd1 )+$signed( { 1'b0,x395 }  )+$signed( { 1'b0,x651 }  )+$signed( -{ 2'b0,x154 }<<<3'd1 )+$signed( { 1'b0,x410 }  )+$signed( { 1'b0,x666 }  )+$signed( -{ 1'b0,x155 } )+$signed(11'd64);
assign y485=temp_y[485][11] ==1'b1 ? 5'd0 :  
        temp_y[485][8] ==1'b1 ? 5'd31 : 
        temp_y[485][2]==1'b1 ? temp_y[485][7:3]+1'b1 : temp_y[485][7:3];
assign temp_y[549] = 
+$signed( -{ 2'b0,x138 }<<<3'd1 )+$signed( -{ 1'b0,x394 } )+$signed( -{ 3'b0,x139 }<<<3'd2)+$signed( { 1'b0,x154 }  )+$signed( { 1'b0,x410 }  )+$signed( { 3'b0,x155 }<<<3'd2 )+$signed(11'd16);
assign y549=temp_y[549][11] ==1'b1 ? 5'd0 :  
        temp_y[549][8] ==1'b1 ? 5'd31 : 
        temp_y[549][2]==1'b1 ? temp_y[549][7:3]+1'b1 : temp_y[549][7:3];
assign temp_y[613] = 
+$signed( { 2'b0,x394 } <<<3'd1 )+$signed( { 2'b0,x650 } <<<3'd1 )+$signed( -{ 1'b0,x139 } )+$signed( -{ 2'b0,x395 }<<<3'd1 )+$signed( -{ 2'b0,x651 }<<<3'd1 )+$signed( { 2'b0,x410 } <<<3'd1 )+$signed( { 1'b0,x666 }  )+$signed( -{ 2'b0,x411 }<<<3'd1 )-$signed(11'd8);
assign y613=temp_y[613][11] ==1'b1 ? 5'd0 :  
        temp_y[613][8] ==1'b1 ? 5'd31 : 
        temp_y[613][2]==1'b1 ? temp_y[613][7:3]+1'b1 : temp_y[613][7:3];
assign temp_y[38] = 
+$signed( -{ 2'b0,x396 }<<<3'd1 )+$signed( -{ 1'b0,x652 } )+$signed( { 1'b0,x141 }  )+$signed( { 1'b0,x397 }  )+$signed( { 1'b0,x653 }  )+$signed( -{ 2'b0,x412 }<<<3'd1 )+$signed( -{ 2'b0,x668 }<<<3'd1 )+$signed( { 2'b0,x413 } <<<3'd1 )+$signed( { 2'b0,x669 } <<<3'd1 )-$signed(11'd16);
assign y38=temp_y[38][11] ==1'b1 ? 5'd0 :  
        temp_y[38][8] ==1'b1 ? 5'd31 : 
        temp_y[38][2]==1'b1 ? temp_y[38][7:3]+1'b1 : temp_y[38][7:3];
assign temp_y[102] = 
+$signed( { 3'b0,x140 }<<<3'd2 )+$signed( -{ 2'b0,x396 }<<<3'd1 )+$signed( -{ 2'b0,x652 }<<<3'd1 )+$signed( { 2'b0,x141 } <<<3'd1 )+$signed( -{ 3'b0,x397 }<<<3'd2)+$signed( { 1'b0,x653 }  )+$signed( -{ 1'b0,x156 } )+$signed( { 1'b0,x668 }  )+$signed( -{ 2'b0,x157 }<<<3'd1 )+$signed( -{ 1'b0,x413 } )+$signed( { 2'b0,x669 } <<<3'd1 )+$signed(11'd24);
assign y102=temp_y[102][11] ==1'b1 ? 5'd0 :  
        temp_y[102][8] ==1'b1 ? 5'd31 : 
        temp_y[102][2]==1'b1 ? temp_y[102][7:3]+1'b1 : temp_y[102][7:3];
assign temp_y[166] = 
+$signed( { 2'b0,x140 } <<<3'd1 )+$signed( { 2'b0,x396 } <<<3'd1 )+$signed( { 1'b0,x652 }  )+$signed( { 2'b0,x141 } <<<3'd1 )+$signed( -{ 1'b0,x397 } )+$signed( { 1'b0,x653 }  )+$signed( -{ 2'b0,x156 }<<<3'd1 )+$signed( -{ 2'b0,x412 }<<<3'd1 )+$signed( -{ 1'b0,x668 } )+$signed( -{ 1'b0,x157 } )+$signed( -{ 1'b0,x413 } )+$signed( -{ 1'b0,x669 } )+$signed(11'd16);
assign y166=temp_y[166][11] ==1'b1 ? 5'd0 :  
        temp_y[166][8] ==1'b1 ? 5'd31 : 
        temp_y[166][2]==1'b1 ? temp_y[166][7:3]+1'b1 : temp_y[166][7:3];
assign temp_y[230] = 
+$signed( { 1'b0,x140 }  )+$signed( -{ 1'b0,x396 } )+$signed( { 1'b0,x141 }  )+$signed( -{ 1'b0,x397 } )+$signed( { 2'b0,x156 } <<<3'd1 )+$signed( -{ 1'b0,x412 } )+$signed( -{ 1'b0,x668 } )+$signed( { 2'b0,x157 } <<<3'd1 )+$signed( -{ 1'b0,x413 } )+$signed( -{ 2'b0,x669 }<<<3'd1 )+$signed(11'd40);
assign y230=temp_y[230][11] ==1'b1 ? 5'd0 :  
        temp_y[230][8] ==1'b1 ? 5'd31 : 
        temp_y[230][2]==1'b1 ? temp_y[230][7:3]+1'b1 : temp_y[230][7:3];
assign temp_y[294] = 
+$signed( -{ 1'b0,x140 } )+$signed( { 2'b0,x396 } <<<3'd1 )+$signed( -{ 1'b0,x652 } )+$signed( -{ 1'b0,x141 } )+$signed( { 2'b0,x397 } <<<3'd1 )+$signed( -{ 2'b0,x653 }<<<3'd1 )+$signed( -{ 1'b0,x156 } )+$signed( { 2'b0,x412 } <<<3'd1 )+$signed( -{ 1'b0,x668 } )+$signed( -{ 2'b0,x157 }<<<3'd1 )+$signed( { 3'b0,x413 }<<<3'd2 )+$signed( -{ 2'b0,x669 }<<<3'd1 )+$signed(11'd32);
assign y294=temp_y[294][11] ==1'b1 ? 5'd0 :  
        temp_y[294][8] ==1'b1 ? 5'd31 : 
        temp_y[294][2]==1'b1 ? temp_y[294][7:3]+1'b1 : temp_y[294][7:3];
assign temp_y[358] = 
+$signed( -{ 1'b0,x140 } )+$signed( -{ 2'b0,x396 }<<<3'd1 )+$signed( -{ 1'b0,x652 } )+$signed( { 1'b0,x141 }  )+$signed( { 2'b0,x397 } <<<3'd1 )+$signed( { 1'b0,x653 }  )+$signed( { 1'b0,x156 }  )+$signed( { 2'b0,x412 } <<<3'd1 )+$signed( { 2'b0,x668 } <<<3'd1 )+$signed( -{ 1'b0,x157 } )+$signed( -{ 2'b0,x413 }<<<3'd1 )+$signed( -{ 1'b0,x669 } )-$signed(11'd68);
assign y358=temp_y[358][11] ==1'b1 ? 5'd0 :  
        temp_y[358][8] ==1'b1 ? 5'd31 : 
        temp_y[358][2]==1'b1 ? temp_y[358][7:3]+1'b1 : temp_y[358][7:3];
assign temp_y[422] = 
+$signed( { 1'b0,x396 }  )+$signed( { 1'b0,x653 }  )+$signed( { 1'b0,x669 }  )-$signed(11'd108);
assign y422=temp_y[422][11] ==1'b1 ? 5'd0 :  
        temp_y[422][8] ==1'b1 ? 5'd31 : 
        temp_y[422][2]==1'b1 ? temp_y[422][7:3]+1'b1 : temp_y[422][7:3];
assign temp_y[486] = 
+$signed( -{ 2'b0,x140 }<<<3'd1 )+$signed( { 2'b0,x652 } <<<3'd1 )+$signed( -{ 2'b0,x141 }<<<3'd1 )+$signed( { 1'b0,x397 }  )+$signed( { 1'b0,x653 }  )+$signed( -{ 2'b0,x156 }<<<3'd1 )+$signed( { 1'b0,x412 }  )+$signed( { 1'b0,x668 }  )+$signed( -{ 1'b0,x157 } )+$signed(11'd64);
assign y486=temp_y[486][11] ==1'b1 ? 5'd0 :  
        temp_y[486][8] ==1'b1 ? 5'd31 : 
        temp_y[486][2]==1'b1 ? temp_y[486][7:3]+1'b1 : temp_y[486][7:3];
assign temp_y[550] = 
+$signed( -{ 2'b0,x140 }<<<3'd1 )+$signed( -{ 1'b0,x396 } )+$signed( -{ 3'b0,x141 }<<<3'd2)+$signed( { 1'b0,x156 }  )+$signed( { 1'b0,x412 }  )+$signed( { 3'b0,x157 }<<<3'd2 )+$signed(11'd16);
assign y550=temp_y[550][11] ==1'b1 ? 5'd0 :  
        temp_y[550][8] ==1'b1 ? 5'd31 : 
        temp_y[550][2]==1'b1 ? temp_y[550][7:3]+1'b1 : temp_y[550][7:3];
assign temp_y[614] = 
+$signed( { 2'b0,x396 } <<<3'd1 )+$signed( { 2'b0,x652 } <<<3'd1 )+$signed( -{ 1'b0,x141 } )+$signed( -{ 2'b0,x397 }<<<3'd1 )+$signed( -{ 2'b0,x653 }<<<3'd1 )+$signed( { 2'b0,x412 } <<<3'd1 )+$signed( { 1'b0,x668 }  )+$signed( -{ 2'b0,x413 }<<<3'd1 )-$signed(11'd8);
assign y614=temp_y[614][11] ==1'b1 ? 5'd0 :  
        temp_y[614][8] ==1'b1 ? 5'd31 : 
        temp_y[614][2]==1'b1 ? temp_y[614][7:3]+1'b1 : temp_y[614][7:3];
assign temp_y[39] = 
+$signed( -{ 2'b0,x398 }<<<3'd1 )+$signed( -{ 1'b0,x654 } )+$signed( { 1'b0,x143 }  )+$signed( { 1'b0,x399 }  )+$signed( { 1'b0,x655 }  )+$signed( -{ 2'b0,x414 }<<<3'd1 )+$signed( -{ 2'b0,x670 }<<<3'd1 )+$signed( { 2'b0,x415 } <<<3'd1 )+$signed( { 2'b0,x671 } <<<3'd1 )-$signed(11'd16);
assign y39=temp_y[39][11] ==1'b1 ? 5'd0 :  
        temp_y[39][8] ==1'b1 ? 5'd31 : 
        temp_y[39][2]==1'b1 ? temp_y[39][7:3]+1'b1 : temp_y[39][7:3];
assign temp_y[103] = 
+$signed( { 3'b0,x142 }<<<3'd2 )+$signed( -{ 2'b0,x398 }<<<3'd1 )+$signed( -{ 2'b0,x654 }<<<3'd1 )+$signed( { 2'b0,x143 } <<<3'd1 )+$signed( -{ 3'b0,x399 }<<<3'd2)+$signed( { 1'b0,x655 }  )+$signed( -{ 1'b0,x158 } )+$signed( { 1'b0,x670 }  )+$signed( -{ 2'b0,x159 }<<<3'd1 )+$signed( -{ 1'b0,x415 } )+$signed( { 2'b0,x671 } <<<3'd1 )+$signed(11'd24);
assign y103=temp_y[103][11] ==1'b1 ? 5'd0 :  
        temp_y[103][8] ==1'b1 ? 5'd31 : 
        temp_y[103][2]==1'b1 ? temp_y[103][7:3]+1'b1 : temp_y[103][7:3];
assign temp_y[167] = 
+$signed( { 2'b0,x142 } <<<3'd1 )+$signed( { 2'b0,x398 } <<<3'd1 )+$signed( { 1'b0,x654 }  )+$signed( { 2'b0,x143 } <<<3'd1 )+$signed( -{ 1'b0,x399 } )+$signed( { 1'b0,x655 }  )+$signed( -{ 2'b0,x158 }<<<3'd1 )+$signed( -{ 2'b0,x414 }<<<3'd1 )+$signed( -{ 1'b0,x670 } )+$signed( -{ 1'b0,x159 } )+$signed( -{ 1'b0,x415 } )+$signed( -{ 1'b0,x671 } )+$signed(11'd16);
assign y167=temp_y[167][11] ==1'b1 ? 5'd0 :  
        temp_y[167][8] ==1'b1 ? 5'd31 : 
        temp_y[167][2]==1'b1 ? temp_y[167][7:3]+1'b1 : temp_y[167][7:3];
assign temp_y[231] = 
+$signed( { 1'b0,x142 }  )+$signed( -{ 1'b0,x398 } )+$signed( { 1'b0,x143 }  )+$signed( -{ 1'b0,x399 } )+$signed( { 2'b0,x158 } <<<3'd1 )+$signed( -{ 1'b0,x414 } )+$signed( -{ 1'b0,x670 } )+$signed( { 2'b0,x159 } <<<3'd1 )+$signed( -{ 1'b0,x415 } )+$signed( -{ 2'b0,x671 }<<<3'd1 )+$signed(11'd40);
assign y231=temp_y[231][11] ==1'b1 ? 5'd0 :  
        temp_y[231][8] ==1'b1 ? 5'd31 : 
        temp_y[231][2]==1'b1 ? temp_y[231][7:3]+1'b1 : temp_y[231][7:3];
assign temp_y[295] = 
+$signed( -{ 1'b0,x142 } )+$signed( { 2'b0,x398 } <<<3'd1 )+$signed( -{ 1'b0,x654 } )+$signed( -{ 1'b0,x143 } )+$signed( { 2'b0,x399 } <<<3'd1 )+$signed( -{ 2'b0,x655 }<<<3'd1 )+$signed( -{ 1'b0,x158 } )+$signed( { 2'b0,x414 } <<<3'd1 )+$signed( -{ 1'b0,x670 } )+$signed( -{ 2'b0,x159 }<<<3'd1 )+$signed( { 3'b0,x415 }<<<3'd2 )+$signed( -{ 2'b0,x671 }<<<3'd1 )+$signed(11'd32);
assign y295=temp_y[295][11] ==1'b1 ? 5'd0 :  
        temp_y[295][8] ==1'b1 ? 5'd31 : 
        temp_y[295][2]==1'b1 ? temp_y[295][7:3]+1'b1 : temp_y[295][7:3];
assign temp_y[359] = 
+$signed( -{ 1'b0,x142 } )+$signed( -{ 2'b0,x398 }<<<3'd1 )+$signed( -{ 1'b0,x654 } )+$signed( { 1'b0,x143 }  )+$signed( { 2'b0,x399 } <<<3'd1 )+$signed( { 1'b0,x655 }  )+$signed( { 1'b0,x158 }  )+$signed( { 2'b0,x414 } <<<3'd1 )+$signed( { 2'b0,x670 } <<<3'd1 )+$signed( -{ 1'b0,x159 } )+$signed( -{ 2'b0,x415 }<<<3'd1 )+$signed( -{ 1'b0,x671 } )-$signed(11'd68);
assign y359=temp_y[359][11] ==1'b1 ? 5'd0 :  
        temp_y[359][8] ==1'b1 ? 5'd31 : 
        temp_y[359][2]==1'b1 ? temp_y[359][7:3]+1'b1 : temp_y[359][7:3];
assign temp_y[423] = 
+$signed( { 1'b0,x398 }  )+$signed( { 1'b0,x655 }  )+$signed( { 1'b0,x671 }  )-$signed(11'd108);
assign y423=temp_y[423][11] ==1'b1 ? 5'd0 :  
        temp_y[423][8] ==1'b1 ? 5'd31 : 
        temp_y[423][2]==1'b1 ? temp_y[423][7:3]+1'b1 : temp_y[423][7:3];
assign temp_y[487] = 
+$signed( -{ 2'b0,x142 }<<<3'd1 )+$signed( { 2'b0,x654 } <<<3'd1 )+$signed( -{ 2'b0,x143 }<<<3'd1 )+$signed( { 1'b0,x399 }  )+$signed( { 1'b0,x655 }  )+$signed( -{ 2'b0,x158 }<<<3'd1 )+$signed( { 1'b0,x414 }  )+$signed( { 1'b0,x670 }  )+$signed( -{ 1'b0,x159 } )+$signed(11'd64);
assign y487=temp_y[487][11] ==1'b1 ? 5'd0 :  
        temp_y[487][8] ==1'b1 ? 5'd31 : 
        temp_y[487][2]==1'b1 ? temp_y[487][7:3]+1'b1 : temp_y[487][7:3];
assign temp_y[551] = 
+$signed( -{ 2'b0,x142 }<<<3'd1 )+$signed( -{ 1'b0,x398 } )+$signed( -{ 3'b0,x143 }<<<3'd2)+$signed( { 1'b0,x158 }  )+$signed( { 1'b0,x414 }  )+$signed( { 3'b0,x159 }<<<3'd2 )+$signed(11'd16);
assign y551=temp_y[551][11] ==1'b1 ? 5'd0 :  
        temp_y[551][8] ==1'b1 ? 5'd31 : 
        temp_y[551][2]==1'b1 ? temp_y[551][7:3]+1'b1 : temp_y[551][7:3];
assign temp_y[615] = 
+$signed( { 2'b0,x398 } <<<3'd1 )+$signed( { 2'b0,x654 } <<<3'd1 )+$signed( -{ 1'b0,x143 } )+$signed( -{ 2'b0,x399 }<<<3'd1 )+$signed( -{ 2'b0,x655 }<<<3'd1 )+$signed( { 2'b0,x414 } <<<3'd1 )+$signed( { 1'b0,x670 }  )+$signed( -{ 2'b0,x415 }<<<3'd1 )-$signed(11'd8);
assign y615=temp_y[615][11] ==1'b1 ? 5'd0 :  
        temp_y[615][8] ==1'b1 ? 5'd31 : 
        temp_y[615][2]==1'b1 ? temp_y[615][7:3]+1'b1 : temp_y[615][7:3];
assign temp_y[40] = 
+$signed( -{ 2'b0,x416 }<<<3'd1 )+$signed( -{ 1'b0,x672 } )+$signed( { 1'b0,x161 }  )+$signed( { 1'b0,x417 }  )+$signed( { 1'b0,x673 }  )+$signed( -{ 2'b0,x432 }<<<3'd1 )+$signed( -{ 2'b0,x688 }<<<3'd1 )+$signed( { 2'b0,x433 } <<<3'd1 )+$signed( { 2'b0,x689 } <<<3'd1 )-$signed(11'd16);
assign y40=temp_y[40][11] ==1'b1 ? 5'd0 :  
        temp_y[40][8] ==1'b1 ? 5'd31 : 
        temp_y[40][2]==1'b1 ? temp_y[40][7:3]+1'b1 : temp_y[40][7:3];
assign temp_y[104] = 
+$signed( { 3'b0,x160 }<<<3'd2 )+$signed( -{ 2'b0,x416 }<<<3'd1 )+$signed( -{ 2'b0,x672 }<<<3'd1 )+$signed( { 2'b0,x161 } <<<3'd1 )+$signed( -{ 3'b0,x417 }<<<3'd2)+$signed( { 1'b0,x673 }  )+$signed( -{ 1'b0,x176 } )+$signed( { 1'b0,x688 }  )+$signed( -{ 2'b0,x177 }<<<3'd1 )+$signed( -{ 1'b0,x433 } )+$signed( { 2'b0,x689 } <<<3'd1 )+$signed(11'd24);
assign y104=temp_y[104][11] ==1'b1 ? 5'd0 :  
        temp_y[104][8] ==1'b1 ? 5'd31 : 
        temp_y[104][2]==1'b1 ? temp_y[104][7:3]+1'b1 : temp_y[104][7:3];
assign temp_y[168] = 
+$signed( { 2'b0,x160 } <<<3'd1 )+$signed( { 2'b0,x416 } <<<3'd1 )+$signed( { 1'b0,x672 }  )+$signed( { 2'b0,x161 } <<<3'd1 )+$signed( -{ 1'b0,x417 } )+$signed( { 1'b0,x673 }  )+$signed( -{ 2'b0,x176 }<<<3'd1 )+$signed( -{ 2'b0,x432 }<<<3'd1 )+$signed( -{ 1'b0,x688 } )+$signed( -{ 1'b0,x177 } )+$signed( -{ 1'b0,x433 } )+$signed( -{ 1'b0,x689 } )+$signed(11'd16);
assign y168=temp_y[168][11] ==1'b1 ? 5'd0 :  
        temp_y[168][8] ==1'b1 ? 5'd31 : 
        temp_y[168][2]==1'b1 ? temp_y[168][7:3]+1'b1 : temp_y[168][7:3];
assign temp_y[232] = 
+$signed( { 1'b0,x160 }  )+$signed( -{ 1'b0,x416 } )+$signed( { 1'b0,x161 }  )+$signed( -{ 1'b0,x417 } )+$signed( { 2'b0,x176 } <<<3'd1 )+$signed( -{ 1'b0,x432 } )+$signed( -{ 1'b0,x688 } )+$signed( { 2'b0,x177 } <<<3'd1 )+$signed( -{ 1'b0,x433 } )+$signed( -{ 2'b0,x689 }<<<3'd1 )+$signed(11'd40);
assign y232=temp_y[232][11] ==1'b1 ? 5'd0 :  
        temp_y[232][8] ==1'b1 ? 5'd31 : 
        temp_y[232][2]==1'b1 ? temp_y[232][7:3]+1'b1 : temp_y[232][7:3];
assign temp_y[296] = 
+$signed( -{ 1'b0,x160 } )+$signed( { 2'b0,x416 } <<<3'd1 )+$signed( -{ 1'b0,x672 } )+$signed( -{ 1'b0,x161 } )+$signed( { 2'b0,x417 } <<<3'd1 )+$signed( -{ 2'b0,x673 }<<<3'd1 )+$signed( -{ 1'b0,x176 } )+$signed( { 2'b0,x432 } <<<3'd1 )+$signed( -{ 1'b0,x688 } )+$signed( -{ 2'b0,x177 }<<<3'd1 )+$signed( { 3'b0,x433 }<<<3'd2 )+$signed( -{ 2'b0,x689 }<<<3'd1 )+$signed(11'd32);
assign y296=temp_y[296][11] ==1'b1 ? 5'd0 :  
        temp_y[296][8] ==1'b1 ? 5'd31 : 
        temp_y[296][2]==1'b1 ? temp_y[296][7:3]+1'b1 : temp_y[296][7:3];
assign temp_y[360] = 
+$signed( -{ 1'b0,x160 } )+$signed( -{ 2'b0,x416 }<<<3'd1 )+$signed( -{ 1'b0,x672 } )+$signed( { 1'b0,x161 }  )+$signed( { 2'b0,x417 } <<<3'd1 )+$signed( { 1'b0,x673 }  )+$signed( { 1'b0,x176 }  )+$signed( { 2'b0,x432 } <<<3'd1 )+$signed( { 2'b0,x688 } <<<3'd1 )+$signed( -{ 1'b0,x177 } )+$signed( -{ 2'b0,x433 }<<<3'd1 )+$signed( -{ 1'b0,x689 } )-$signed(11'd68);
assign y360=temp_y[360][11] ==1'b1 ? 5'd0 :  
        temp_y[360][8] ==1'b1 ? 5'd31 : 
        temp_y[360][2]==1'b1 ? temp_y[360][7:3]+1'b1 : temp_y[360][7:3];
assign temp_y[424] = 
+$signed( { 1'b0,x416 }  )+$signed( { 1'b0,x673 }  )+$signed( { 1'b0,x689 }  )-$signed(11'd108);
assign y424=temp_y[424][11] ==1'b1 ? 5'd0 :  
        temp_y[424][8] ==1'b1 ? 5'd31 : 
        temp_y[424][2]==1'b1 ? temp_y[424][7:3]+1'b1 : temp_y[424][7:3];
assign temp_y[488] = 
+$signed( -{ 2'b0,x160 }<<<3'd1 )+$signed( { 2'b0,x672 } <<<3'd1 )+$signed( -{ 2'b0,x161 }<<<3'd1 )+$signed( { 1'b0,x417 }  )+$signed( { 1'b0,x673 }  )+$signed( -{ 2'b0,x176 }<<<3'd1 )+$signed( { 1'b0,x432 }  )+$signed( { 1'b0,x688 }  )+$signed( -{ 1'b0,x177 } )+$signed(11'd64);
assign y488=temp_y[488][11] ==1'b1 ? 5'd0 :  
        temp_y[488][8] ==1'b1 ? 5'd31 : 
        temp_y[488][2]==1'b1 ? temp_y[488][7:3]+1'b1 : temp_y[488][7:3];
assign temp_y[552] = 
+$signed( -{ 2'b0,x160 }<<<3'd1 )+$signed( -{ 1'b0,x416 } )+$signed( -{ 3'b0,x161 }<<<3'd2)+$signed( { 1'b0,x176 }  )+$signed( { 1'b0,x432 }  )+$signed( { 3'b0,x177 }<<<3'd2 )+$signed(11'd16);
assign y552=temp_y[552][11] ==1'b1 ? 5'd0 :  
        temp_y[552][8] ==1'b1 ? 5'd31 : 
        temp_y[552][2]==1'b1 ? temp_y[552][7:3]+1'b1 : temp_y[552][7:3];
assign temp_y[616] = 
+$signed( { 2'b0,x416 } <<<3'd1 )+$signed( { 2'b0,x672 } <<<3'd1 )+$signed( -{ 1'b0,x161 } )+$signed( -{ 2'b0,x417 }<<<3'd1 )+$signed( -{ 2'b0,x673 }<<<3'd1 )+$signed( { 2'b0,x432 } <<<3'd1 )+$signed( { 1'b0,x688 }  )+$signed( -{ 2'b0,x433 }<<<3'd1 )-$signed(11'd8);
assign y616=temp_y[616][11] ==1'b1 ? 5'd0 :  
        temp_y[616][8] ==1'b1 ? 5'd31 : 
        temp_y[616][2]==1'b1 ? temp_y[616][7:3]+1'b1 : temp_y[616][7:3];
assign temp_y[41] = 
+$signed( -{ 2'b0,x418 }<<<3'd1 )+$signed( -{ 1'b0,x674 } )+$signed( { 1'b0,x163 }  )+$signed( { 1'b0,x419 }  )+$signed( { 1'b0,x675 }  )+$signed( -{ 2'b0,x434 }<<<3'd1 )+$signed( -{ 2'b0,x690 }<<<3'd1 )+$signed( { 2'b0,x435 } <<<3'd1 )+$signed( { 2'b0,x691 } <<<3'd1 )-$signed(11'd16);
assign y41=temp_y[41][11] ==1'b1 ? 5'd0 :  
        temp_y[41][8] ==1'b1 ? 5'd31 : 
        temp_y[41][2]==1'b1 ? temp_y[41][7:3]+1'b1 : temp_y[41][7:3];
assign temp_y[105] = 
+$signed( { 3'b0,x162 }<<<3'd2 )+$signed( -{ 2'b0,x418 }<<<3'd1 )+$signed( -{ 2'b0,x674 }<<<3'd1 )+$signed( { 2'b0,x163 } <<<3'd1 )+$signed( -{ 3'b0,x419 }<<<3'd2)+$signed( { 1'b0,x675 }  )+$signed( -{ 1'b0,x178 } )+$signed( { 1'b0,x690 }  )+$signed( -{ 2'b0,x179 }<<<3'd1 )+$signed( -{ 1'b0,x435 } )+$signed( { 2'b0,x691 } <<<3'd1 )+$signed(11'd24);
assign y105=temp_y[105][11] ==1'b1 ? 5'd0 :  
        temp_y[105][8] ==1'b1 ? 5'd31 : 
        temp_y[105][2]==1'b1 ? temp_y[105][7:3]+1'b1 : temp_y[105][7:3];
assign temp_y[169] = 
+$signed( { 2'b0,x162 } <<<3'd1 )+$signed( { 2'b0,x418 } <<<3'd1 )+$signed( { 1'b0,x674 }  )+$signed( { 2'b0,x163 } <<<3'd1 )+$signed( -{ 1'b0,x419 } )+$signed( { 1'b0,x675 }  )+$signed( -{ 2'b0,x178 }<<<3'd1 )+$signed( -{ 2'b0,x434 }<<<3'd1 )+$signed( -{ 1'b0,x690 } )+$signed( -{ 1'b0,x179 } )+$signed( -{ 1'b0,x435 } )+$signed( -{ 1'b0,x691 } )+$signed(11'd16);
assign y169=temp_y[169][11] ==1'b1 ? 5'd0 :  
        temp_y[169][8] ==1'b1 ? 5'd31 : 
        temp_y[169][2]==1'b1 ? temp_y[169][7:3]+1'b1 : temp_y[169][7:3];
assign temp_y[233] = 
+$signed( { 1'b0,x162 }  )+$signed( -{ 1'b0,x418 } )+$signed( { 1'b0,x163 }  )+$signed( -{ 1'b0,x419 } )+$signed( { 2'b0,x178 } <<<3'd1 )+$signed( -{ 1'b0,x434 } )+$signed( -{ 1'b0,x690 } )+$signed( { 2'b0,x179 } <<<3'd1 )+$signed( -{ 1'b0,x435 } )+$signed( -{ 2'b0,x691 }<<<3'd1 )+$signed(11'd40);
assign y233=temp_y[233][11] ==1'b1 ? 5'd0 :  
        temp_y[233][8] ==1'b1 ? 5'd31 : 
        temp_y[233][2]==1'b1 ? temp_y[233][7:3]+1'b1 : temp_y[233][7:3];
assign temp_y[297] = 
+$signed( -{ 1'b0,x162 } )+$signed( { 2'b0,x418 } <<<3'd1 )+$signed( -{ 1'b0,x674 } )+$signed( -{ 1'b0,x163 } )+$signed( { 2'b0,x419 } <<<3'd1 )+$signed( -{ 2'b0,x675 }<<<3'd1 )+$signed( -{ 1'b0,x178 } )+$signed( { 2'b0,x434 } <<<3'd1 )+$signed( -{ 1'b0,x690 } )+$signed( -{ 2'b0,x179 }<<<3'd1 )+$signed( { 3'b0,x435 }<<<3'd2 )+$signed( -{ 2'b0,x691 }<<<3'd1 )+$signed(11'd32);
assign y297=temp_y[297][11] ==1'b1 ? 5'd0 :  
        temp_y[297][8] ==1'b1 ? 5'd31 : 
        temp_y[297][2]==1'b1 ? temp_y[297][7:3]+1'b1 : temp_y[297][7:3];
assign temp_y[361] = 
+$signed( -{ 1'b0,x162 } )+$signed( -{ 2'b0,x418 }<<<3'd1 )+$signed( -{ 1'b0,x674 } )+$signed( { 1'b0,x163 }  )+$signed( { 2'b0,x419 } <<<3'd1 )+$signed( { 1'b0,x675 }  )+$signed( { 1'b0,x178 }  )+$signed( { 2'b0,x434 } <<<3'd1 )+$signed( { 2'b0,x690 } <<<3'd1 )+$signed( -{ 1'b0,x179 } )+$signed( -{ 2'b0,x435 }<<<3'd1 )+$signed( -{ 1'b0,x691 } )-$signed(11'd68);
assign y361=temp_y[361][11] ==1'b1 ? 5'd0 :  
        temp_y[361][8] ==1'b1 ? 5'd31 : 
        temp_y[361][2]==1'b1 ? temp_y[361][7:3]+1'b1 : temp_y[361][7:3];
assign temp_y[425] = 
+$signed( { 1'b0,x418 }  )+$signed( { 1'b0,x675 }  )+$signed( { 1'b0,x691 }  )-$signed(11'd108);
assign y425=temp_y[425][11] ==1'b1 ? 5'd0 :  
        temp_y[425][8] ==1'b1 ? 5'd31 : 
        temp_y[425][2]==1'b1 ? temp_y[425][7:3]+1'b1 : temp_y[425][7:3];
assign temp_y[489] = 
+$signed( -{ 2'b0,x162 }<<<3'd1 )+$signed( { 2'b0,x674 } <<<3'd1 )+$signed( -{ 2'b0,x163 }<<<3'd1 )+$signed( { 1'b0,x419 }  )+$signed( { 1'b0,x675 }  )+$signed( -{ 2'b0,x178 }<<<3'd1 )+$signed( { 1'b0,x434 }  )+$signed( { 1'b0,x690 }  )+$signed( -{ 1'b0,x179 } )+$signed(11'd64);
assign y489=temp_y[489][11] ==1'b1 ? 5'd0 :  
        temp_y[489][8] ==1'b1 ? 5'd31 : 
        temp_y[489][2]==1'b1 ? temp_y[489][7:3]+1'b1 : temp_y[489][7:3];
assign temp_y[553] = 
+$signed( -{ 2'b0,x162 }<<<3'd1 )+$signed( -{ 1'b0,x418 } )+$signed( -{ 3'b0,x163 }<<<3'd2)+$signed( { 1'b0,x178 }  )+$signed( { 1'b0,x434 }  )+$signed( { 3'b0,x179 }<<<3'd2 )+$signed(11'd16);
assign y553=temp_y[553][11] ==1'b1 ? 5'd0 :  
        temp_y[553][8] ==1'b1 ? 5'd31 : 
        temp_y[553][2]==1'b1 ? temp_y[553][7:3]+1'b1 : temp_y[553][7:3];
assign temp_y[617] = 
+$signed( { 2'b0,x418 } <<<3'd1 )+$signed( { 2'b0,x674 } <<<3'd1 )+$signed( -{ 1'b0,x163 } )+$signed( -{ 2'b0,x419 }<<<3'd1 )+$signed( -{ 2'b0,x675 }<<<3'd1 )+$signed( { 2'b0,x434 } <<<3'd1 )+$signed( { 1'b0,x690 }  )+$signed( -{ 2'b0,x435 }<<<3'd1 )-$signed(11'd8);
assign y617=temp_y[617][11] ==1'b1 ? 5'd0 :  
        temp_y[617][8] ==1'b1 ? 5'd31 : 
        temp_y[617][2]==1'b1 ? temp_y[617][7:3]+1'b1 : temp_y[617][7:3];
assign temp_y[42] = 
+$signed( -{ 2'b0,x420 }<<<3'd1 )+$signed( -{ 1'b0,x676 } )+$signed( { 1'b0,x165 }  )+$signed( { 1'b0,x421 }  )+$signed( { 1'b0,x677 }  )+$signed( -{ 2'b0,x436 }<<<3'd1 )+$signed( -{ 2'b0,x692 }<<<3'd1 )+$signed( { 2'b0,x437 } <<<3'd1 )+$signed( { 2'b0,x693 } <<<3'd1 )-$signed(11'd16);
assign y42=temp_y[42][11] ==1'b1 ? 5'd0 :  
        temp_y[42][8] ==1'b1 ? 5'd31 : 
        temp_y[42][2]==1'b1 ? temp_y[42][7:3]+1'b1 : temp_y[42][7:3];
assign temp_y[106] = 
+$signed( { 3'b0,x164 }<<<3'd2 )+$signed( -{ 2'b0,x420 }<<<3'd1 )+$signed( -{ 2'b0,x676 }<<<3'd1 )+$signed( { 2'b0,x165 } <<<3'd1 )+$signed( -{ 3'b0,x421 }<<<3'd2)+$signed( { 1'b0,x677 }  )+$signed( -{ 1'b0,x180 } )+$signed( { 1'b0,x692 }  )+$signed( -{ 2'b0,x181 }<<<3'd1 )+$signed( -{ 1'b0,x437 } )+$signed( { 2'b0,x693 } <<<3'd1 )+$signed(11'd24);
assign y106=temp_y[106][11] ==1'b1 ? 5'd0 :  
        temp_y[106][8] ==1'b1 ? 5'd31 : 
        temp_y[106][2]==1'b1 ? temp_y[106][7:3]+1'b1 : temp_y[106][7:3];
assign temp_y[170] = 
+$signed( { 2'b0,x164 } <<<3'd1 )+$signed( { 2'b0,x420 } <<<3'd1 )+$signed( { 1'b0,x676 }  )+$signed( { 2'b0,x165 } <<<3'd1 )+$signed( -{ 1'b0,x421 } )+$signed( { 1'b0,x677 }  )+$signed( -{ 2'b0,x180 }<<<3'd1 )+$signed( -{ 2'b0,x436 }<<<3'd1 )+$signed( -{ 1'b0,x692 } )+$signed( -{ 1'b0,x181 } )+$signed( -{ 1'b0,x437 } )+$signed( -{ 1'b0,x693 } )+$signed(11'd16);
assign y170=temp_y[170][11] ==1'b1 ? 5'd0 :  
        temp_y[170][8] ==1'b1 ? 5'd31 : 
        temp_y[170][2]==1'b1 ? temp_y[170][7:3]+1'b1 : temp_y[170][7:3];
assign temp_y[234] = 
+$signed( { 1'b0,x164 }  )+$signed( -{ 1'b0,x420 } )+$signed( { 1'b0,x165 }  )+$signed( -{ 1'b0,x421 } )+$signed( { 2'b0,x180 } <<<3'd1 )+$signed( -{ 1'b0,x436 } )+$signed( -{ 1'b0,x692 } )+$signed( { 2'b0,x181 } <<<3'd1 )+$signed( -{ 1'b0,x437 } )+$signed( -{ 2'b0,x693 }<<<3'd1 )+$signed(11'd40);
assign y234=temp_y[234][11] ==1'b1 ? 5'd0 :  
        temp_y[234][8] ==1'b1 ? 5'd31 : 
        temp_y[234][2]==1'b1 ? temp_y[234][7:3]+1'b1 : temp_y[234][7:3];
assign temp_y[298] = 
+$signed( -{ 1'b0,x164 } )+$signed( { 2'b0,x420 } <<<3'd1 )+$signed( -{ 1'b0,x676 } )+$signed( -{ 1'b0,x165 } )+$signed( { 2'b0,x421 } <<<3'd1 )+$signed( -{ 2'b0,x677 }<<<3'd1 )+$signed( -{ 1'b0,x180 } )+$signed( { 2'b0,x436 } <<<3'd1 )+$signed( -{ 1'b0,x692 } )+$signed( -{ 2'b0,x181 }<<<3'd1 )+$signed( { 3'b0,x437 }<<<3'd2 )+$signed( -{ 2'b0,x693 }<<<3'd1 )+$signed(11'd32);
assign y298=temp_y[298][11] ==1'b1 ? 5'd0 :  
        temp_y[298][8] ==1'b1 ? 5'd31 : 
        temp_y[298][2]==1'b1 ? temp_y[298][7:3]+1'b1 : temp_y[298][7:3];
assign temp_y[362] = 
+$signed( -{ 1'b0,x164 } )+$signed( -{ 2'b0,x420 }<<<3'd1 )+$signed( -{ 1'b0,x676 } )+$signed( { 1'b0,x165 }  )+$signed( { 2'b0,x421 } <<<3'd1 )+$signed( { 1'b0,x677 }  )+$signed( { 1'b0,x180 }  )+$signed( { 2'b0,x436 } <<<3'd1 )+$signed( { 2'b0,x692 } <<<3'd1 )+$signed( -{ 1'b0,x181 } )+$signed( -{ 2'b0,x437 }<<<3'd1 )+$signed( -{ 1'b0,x693 } )-$signed(11'd68);
assign y362=temp_y[362][11] ==1'b1 ? 5'd0 :  
        temp_y[362][8] ==1'b1 ? 5'd31 : 
        temp_y[362][2]==1'b1 ? temp_y[362][7:3]+1'b1 : temp_y[362][7:3];
assign temp_y[426] = 
+$signed( { 1'b0,x420 }  )+$signed( { 1'b0,x677 }  )+$signed( { 1'b0,x693 }  )-$signed(11'd108);
assign y426=temp_y[426][11] ==1'b1 ? 5'd0 :  
        temp_y[426][8] ==1'b1 ? 5'd31 : 
        temp_y[426][2]==1'b1 ? temp_y[426][7:3]+1'b1 : temp_y[426][7:3];
assign temp_y[490] = 
+$signed( -{ 2'b0,x164 }<<<3'd1 )+$signed( { 2'b0,x676 } <<<3'd1 )+$signed( -{ 2'b0,x165 }<<<3'd1 )+$signed( { 1'b0,x421 }  )+$signed( { 1'b0,x677 }  )+$signed( -{ 2'b0,x180 }<<<3'd1 )+$signed( { 1'b0,x436 }  )+$signed( { 1'b0,x692 }  )+$signed( -{ 1'b0,x181 } )+$signed(11'd64);
assign y490=temp_y[490][11] ==1'b1 ? 5'd0 :  
        temp_y[490][8] ==1'b1 ? 5'd31 : 
        temp_y[490][2]==1'b1 ? temp_y[490][7:3]+1'b1 : temp_y[490][7:3];
assign temp_y[554] = 
+$signed( -{ 2'b0,x164 }<<<3'd1 )+$signed( -{ 1'b0,x420 } )+$signed( -{ 3'b0,x165 }<<<3'd2)+$signed( { 1'b0,x180 }  )+$signed( { 1'b0,x436 }  )+$signed( { 3'b0,x181 }<<<3'd2 )+$signed(11'd16);
assign y554=temp_y[554][11] ==1'b1 ? 5'd0 :  
        temp_y[554][8] ==1'b1 ? 5'd31 : 
        temp_y[554][2]==1'b1 ? temp_y[554][7:3]+1'b1 : temp_y[554][7:3];
assign temp_y[618] = 
+$signed( { 2'b0,x420 } <<<3'd1 )+$signed( { 2'b0,x676 } <<<3'd1 )+$signed( -{ 1'b0,x165 } )+$signed( -{ 2'b0,x421 }<<<3'd1 )+$signed( -{ 2'b0,x677 }<<<3'd1 )+$signed( { 2'b0,x436 } <<<3'd1 )+$signed( { 1'b0,x692 }  )+$signed( -{ 2'b0,x437 }<<<3'd1 )-$signed(11'd8);
assign y618=temp_y[618][11] ==1'b1 ? 5'd0 :  
        temp_y[618][8] ==1'b1 ? 5'd31 : 
        temp_y[618][2]==1'b1 ? temp_y[618][7:3]+1'b1 : temp_y[618][7:3];
assign temp_y[43] = 
+$signed( -{ 2'b0,x422 }<<<3'd1 )+$signed( -{ 1'b0,x678 } )+$signed( { 1'b0,x167 }  )+$signed( { 1'b0,x423 }  )+$signed( { 1'b0,x679 }  )+$signed( -{ 2'b0,x438 }<<<3'd1 )+$signed( -{ 2'b0,x694 }<<<3'd1 )+$signed( { 2'b0,x439 } <<<3'd1 )+$signed( { 2'b0,x695 } <<<3'd1 )-$signed(11'd16);
assign y43=temp_y[43][11] ==1'b1 ? 5'd0 :  
        temp_y[43][8] ==1'b1 ? 5'd31 : 
        temp_y[43][2]==1'b1 ? temp_y[43][7:3]+1'b1 : temp_y[43][7:3];
assign temp_y[107] = 
+$signed( { 3'b0,x166 }<<<3'd2 )+$signed( -{ 2'b0,x422 }<<<3'd1 )+$signed( -{ 2'b0,x678 }<<<3'd1 )+$signed( { 2'b0,x167 } <<<3'd1 )+$signed( -{ 3'b0,x423 }<<<3'd2)+$signed( { 1'b0,x679 }  )+$signed( -{ 1'b0,x182 } )+$signed( { 1'b0,x694 }  )+$signed( -{ 2'b0,x183 }<<<3'd1 )+$signed( -{ 1'b0,x439 } )+$signed( { 2'b0,x695 } <<<3'd1 )+$signed(11'd24);
assign y107=temp_y[107][11] ==1'b1 ? 5'd0 :  
        temp_y[107][8] ==1'b1 ? 5'd31 : 
        temp_y[107][2]==1'b1 ? temp_y[107][7:3]+1'b1 : temp_y[107][7:3];
assign temp_y[171] = 
+$signed( { 2'b0,x166 } <<<3'd1 )+$signed( { 2'b0,x422 } <<<3'd1 )+$signed( { 1'b0,x678 }  )+$signed( { 2'b0,x167 } <<<3'd1 )+$signed( -{ 1'b0,x423 } )+$signed( { 1'b0,x679 }  )+$signed( -{ 2'b0,x182 }<<<3'd1 )+$signed( -{ 2'b0,x438 }<<<3'd1 )+$signed( -{ 1'b0,x694 } )+$signed( -{ 1'b0,x183 } )+$signed( -{ 1'b0,x439 } )+$signed( -{ 1'b0,x695 } )+$signed(11'd16);
assign y171=temp_y[171][11] ==1'b1 ? 5'd0 :  
        temp_y[171][8] ==1'b1 ? 5'd31 : 
        temp_y[171][2]==1'b1 ? temp_y[171][7:3]+1'b1 : temp_y[171][7:3];
assign temp_y[235] = 
+$signed( { 1'b0,x166 }  )+$signed( -{ 1'b0,x422 } )+$signed( { 1'b0,x167 }  )+$signed( -{ 1'b0,x423 } )+$signed( { 2'b0,x182 } <<<3'd1 )+$signed( -{ 1'b0,x438 } )+$signed( -{ 1'b0,x694 } )+$signed( { 2'b0,x183 } <<<3'd1 )+$signed( -{ 1'b0,x439 } )+$signed( -{ 2'b0,x695 }<<<3'd1 )+$signed(11'd40);
assign y235=temp_y[235][11] ==1'b1 ? 5'd0 :  
        temp_y[235][8] ==1'b1 ? 5'd31 : 
        temp_y[235][2]==1'b1 ? temp_y[235][7:3]+1'b1 : temp_y[235][7:3];
assign temp_y[299] = 
+$signed( -{ 1'b0,x166 } )+$signed( { 2'b0,x422 } <<<3'd1 )+$signed( -{ 1'b0,x678 } )+$signed( -{ 1'b0,x167 } )+$signed( { 2'b0,x423 } <<<3'd1 )+$signed( -{ 2'b0,x679 }<<<3'd1 )+$signed( -{ 1'b0,x182 } )+$signed( { 2'b0,x438 } <<<3'd1 )+$signed( -{ 1'b0,x694 } )+$signed( -{ 2'b0,x183 }<<<3'd1 )+$signed( { 3'b0,x439 }<<<3'd2 )+$signed( -{ 2'b0,x695 }<<<3'd1 )+$signed(11'd32);
assign y299=temp_y[299][11] ==1'b1 ? 5'd0 :  
        temp_y[299][8] ==1'b1 ? 5'd31 : 
        temp_y[299][2]==1'b1 ? temp_y[299][7:3]+1'b1 : temp_y[299][7:3];
assign temp_y[363] = 
+$signed( -{ 1'b0,x166 } )+$signed( -{ 2'b0,x422 }<<<3'd1 )+$signed( -{ 1'b0,x678 } )+$signed( { 1'b0,x167 }  )+$signed( { 2'b0,x423 } <<<3'd1 )+$signed( { 1'b0,x679 }  )+$signed( { 1'b0,x182 }  )+$signed( { 2'b0,x438 } <<<3'd1 )+$signed( { 2'b0,x694 } <<<3'd1 )+$signed( -{ 1'b0,x183 } )+$signed( -{ 2'b0,x439 }<<<3'd1 )+$signed( -{ 1'b0,x695 } )-$signed(11'd68);
assign y363=temp_y[363][11] ==1'b1 ? 5'd0 :  
        temp_y[363][8] ==1'b1 ? 5'd31 : 
        temp_y[363][2]==1'b1 ? temp_y[363][7:3]+1'b1 : temp_y[363][7:3];
assign temp_y[427] = 
+$signed( { 1'b0,x422 }  )+$signed( { 1'b0,x679 }  )+$signed( { 1'b0,x695 }  )-$signed(11'd108);
assign y427=temp_y[427][11] ==1'b1 ? 5'd0 :  
        temp_y[427][8] ==1'b1 ? 5'd31 : 
        temp_y[427][2]==1'b1 ? temp_y[427][7:3]+1'b1 : temp_y[427][7:3];
assign temp_y[491] = 
+$signed( -{ 2'b0,x166 }<<<3'd1 )+$signed( { 2'b0,x678 } <<<3'd1 )+$signed( -{ 2'b0,x167 }<<<3'd1 )+$signed( { 1'b0,x423 }  )+$signed( { 1'b0,x679 }  )+$signed( -{ 2'b0,x182 }<<<3'd1 )+$signed( { 1'b0,x438 }  )+$signed( { 1'b0,x694 }  )+$signed( -{ 1'b0,x183 } )+$signed(11'd64);
assign y491=temp_y[491][11] ==1'b1 ? 5'd0 :  
        temp_y[491][8] ==1'b1 ? 5'd31 : 
        temp_y[491][2]==1'b1 ? temp_y[491][7:3]+1'b1 : temp_y[491][7:3];
assign temp_y[555] = 
+$signed( -{ 2'b0,x166 }<<<3'd1 )+$signed( -{ 1'b0,x422 } )+$signed( -{ 3'b0,x167 }<<<3'd2)+$signed( { 1'b0,x182 }  )+$signed( { 1'b0,x438 }  )+$signed( { 3'b0,x183 }<<<3'd2 )+$signed(11'd16);
assign y555=temp_y[555][11] ==1'b1 ? 5'd0 :  
        temp_y[555][8] ==1'b1 ? 5'd31 : 
        temp_y[555][2]==1'b1 ? temp_y[555][7:3]+1'b1 : temp_y[555][7:3];
assign temp_y[619] = 
+$signed( { 2'b0,x422 } <<<3'd1 )+$signed( { 2'b0,x678 } <<<3'd1 )+$signed( -{ 1'b0,x167 } )+$signed( -{ 2'b0,x423 }<<<3'd1 )+$signed( -{ 2'b0,x679 }<<<3'd1 )+$signed( { 2'b0,x438 } <<<3'd1 )+$signed( { 1'b0,x694 }  )+$signed( -{ 2'b0,x439 }<<<3'd1 )-$signed(11'd8);
assign y619=temp_y[619][11] ==1'b1 ? 5'd0 :  
        temp_y[619][8] ==1'b1 ? 5'd31 : 
        temp_y[619][2]==1'b1 ? temp_y[619][7:3]+1'b1 : temp_y[619][7:3];
assign temp_y[44] = 
+$signed( -{ 2'b0,x424 }<<<3'd1 )+$signed( -{ 1'b0,x680 } )+$signed( { 1'b0,x169 }  )+$signed( { 1'b0,x425 }  )+$signed( { 1'b0,x681 }  )+$signed( -{ 2'b0,x440 }<<<3'd1 )+$signed( -{ 2'b0,x696 }<<<3'd1 )+$signed( { 2'b0,x441 } <<<3'd1 )+$signed( { 2'b0,x697 } <<<3'd1 )-$signed(11'd16);
assign y44=temp_y[44][11] ==1'b1 ? 5'd0 :  
        temp_y[44][8] ==1'b1 ? 5'd31 : 
        temp_y[44][2]==1'b1 ? temp_y[44][7:3]+1'b1 : temp_y[44][7:3];
assign temp_y[108] = 
+$signed( { 3'b0,x168 }<<<3'd2 )+$signed( -{ 2'b0,x424 }<<<3'd1 )+$signed( -{ 2'b0,x680 }<<<3'd1 )+$signed( { 2'b0,x169 } <<<3'd1 )+$signed( -{ 3'b0,x425 }<<<3'd2)+$signed( { 1'b0,x681 }  )+$signed( -{ 1'b0,x184 } )+$signed( { 1'b0,x696 }  )+$signed( -{ 2'b0,x185 }<<<3'd1 )+$signed( -{ 1'b0,x441 } )+$signed( { 2'b0,x697 } <<<3'd1 )+$signed(11'd24);
assign y108=temp_y[108][11] ==1'b1 ? 5'd0 :  
        temp_y[108][8] ==1'b1 ? 5'd31 : 
        temp_y[108][2]==1'b1 ? temp_y[108][7:3]+1'b1 : temp_y[108][7:3];
assign temp_y[172] = 
+$signed( { 2'b0,x168 } <<<3'd1 )+$signed( { 2'b0,x424 } <<<3'd1 )+$signed( { 1'b0,x680 }  )+$signed( { 2'b0,x169 } <<<3'd1 )+$signed( -{ 1'b0,x425 } )+$signed( { 1'b0,x681 }  )+$signed( -{ 2'b0,x184 }<<<3'd1 )+$signed( -{ 2'b0,x440 }<<<3'd1 )+$signed( -{ 1'b0,x696 } )+$signed( -{ 1'b0,x185 } )+$signed( -{ 1'b0,x441 } )+$signed( -{ 1'b0,x697 } )+$signed(11'd16);
assign y172=temp_y[172][11] ==1'b1 ? 5'd0 :  
        temp_y[172][8] ==1'b1 ? 5'd31 : 
        temp_y[172][2]==1'b1 ? temp_y[172][7:3]+1'b1 : temp_y[172][7:3];
assign temp_y[236] = 
+$signed( { 1'b0,x168 }  )+$signed( -{ 1'b0,x424 } )+$signed( { 1'b0,x169 }  )+$signed( -{ 1'b0,x425 } )+$signed( { 2'b0,x184 } <<<3'd1 )+$signed( -{ 1'b0,x440 } )+$signed( -{ 1'b0,x696 } )+$signed( { 2'b0,x185 } <<<3'd1 )+$signed( -{ 1'b0,x441 } )+$signed( -{ 2'b0,x697 }<<<3'd1 )+$signed(11'd40);
assign y236=temp_y[236][11] ==1'b1 ? 5'd0 :  
        temp_y[236][8] ==1'b1 ? 5'd31 : 
        temp_y[236][2]==1'b1 ? temp_y[236][7:3]+1'b1 : temp_y[236][7:3];
assign temp_y[300] = 
+$signed( -{ 1'b0,x168 } )+$signed( { 2'b0,x424 } <<<3'd1 )+$signed( -{ 1'b0,x680 } )+$signed( -{ 1'b0,x169 } )+$signed( { 2'b0,x425 } <<<3'd1 )+$signed( -{ 2'b0,x681 }<<<3'd1 )+$signed( -{ 1'b0,x184 } )+$signed( { 2'b0,x440 } <<<3'd1 )+$signed( -{ 1'b0,x696 } )+$signed( -{ 2'b0,x185 }<<<3'd1 )+$signed( { 3'b0,x441 }<<<3'd2 )+$signed( -{ 2'b0,x697 }<<<3'd1 )+$signed(11'd32);
assign y300=temp_y[300][11] ==1'b1 ? 5'd0 :  
        temp_y[300][8] ==1'b1 ? 5'd31 : 
        temp_y[300][2]==1'b1 ? temp_y[300][7:3]+1'b1 : temp_y[300][7:3];
assign temp_y[364] = 
+$signed( -{ 1'b0,x168 } )+$signed( -{ 2'b0,x424 }<<<3'd1 )+$signed( -{ 1'b0,x680 } )+$signed( { 1'b0,x169 }  )+$signed( { 2'b0,x425 } <<<3'd1 )+$signed( { 1'b0,x681 }  )+$signed( { 1'b0,x184 }  )+$signed( { 2'b0,x440 } <<<3'd1 )+$signed( { 2'b0,x696 } <<<3'd1 )+$signed( -{ 1'b0,x185 } )+$signed( -{ 2'b0,x441 }<<<3'd1 )+$signed( -{ 1'b0,x697 } )-$signed(11'd68);
assign y364=temp_y[364][11] ==1'b1 ? 5'd0 :  
        temp_y[364][8] ==1'b1 ? 5'd31 : 
        temp_y[364][2]==1'b1 ? temp_y[364][7:3]+1'b1 : temp_y[364][7:3];
assign temp_y[428] = 
+$signed( { 1'b0,x424 }  )+$signed( { 1'b0,x681 }  )+$signed( { 1'b0,x697 }  )-$signed(11'd108);
assign y428=temp_y[428][11] ==1'b1 ? 5'd0 :  
        temp_y[428][8] ==1'b1 ? 5'd31 : 
        temp_y[428][2]==1'b1 ? temp_y[428][7:3]+1'b1 : temp_y[428][7:3];
assign temp_y[492] = 
+$signed( -{ 2'b0,x168 }<<<3'd1 )+$signed( { 2'b0,x680 } <<<3'd1 )+$signed( -{ 2'b0,x169 }<<<3'd1 )+$signed( { 1'b0,x425 }  )+$signed( { 1'b0,x681 }  )+$signed( -{ 2'b0,x184 }<<<3'd1 )+$signed( { 1'b0,x440 }  )+$signed( { 1'b0,x696 }  )+$signed( -{ 1'b0,x185 } )+$signed(11'd64);
assign y492=temp_y[492][11] ==1'b1 ? 5'd0 :  
        temp_y[492][8] ==1'b1 ? 5'd31 : 
        temp_y[492][2]==1'b1 ? temp_y[492][7:3]+1'b1 : temp_y[492][7:3];
assign temp_y[556] = 
+$signed( -{ 2'b0,x168 }<<<3'd1 )+$signed( -{ 1'b0,x424 } )+$signed( -{ 3'b0,x169 }<<<3'd2)+$signed( { 1'b0,x184 }  )+$signed( { 1'b0,x440 }  )+$signed( { 3'b0,x185 }<<<3'd2 )+$signed(11'd16);
assign y556=temp_y[556][11] ==1'b1 ? 5'd0 :  
        temp_y[556][8] ==1'b1 ? 5'd31 : 
        temp_y[556][2]==1'b1 ? temp_y[556][7:3]+1'b1 : temp_y[556][7:3];
assign temp_y[620] = 
+$signed( { 2'b0,x424 } <<<3'd1 )+$signed( { 2'b0,x680 } <<<3'd1 )+$signed( -{ 1'b0,x169 } )+$signed( -{ 2'b0,x425 }<<<3'd1 )+$signed( -{ 2'b0,x681 }<<<3'd1 )+$signed( { 2'b0,x440 } <<<3'd1 )+$signed( { 1'b0,x696 }  )+$signed( -{ 2'b0,x441 }<<<3'd1 )-$signed(11'd8);
assign y620=temp_y[620][11] ==1'b1 ? 5'd0 :  
        temp_y[620][8] ==1'b1 ? 5'd31 : 
        temp_y[620][2]==1'b1 ? temp_y[620][7:3]+1'b1 : temp_y[620][7:3];
assign temp_y[45] = 
+$signed( -{ 2'b0,x426 }<<<3'd1 )+$signed( -{ 1'b0,x682 } )+$signed( { 1'b0,x171 }  )+$signed( { 1'b0,x427 }  )+$signed( { 1'b0,x683 }  )+$signed( -{ 2'b0,x442 }<<<3'd1 )+$signed( -{ 2'b0,x698 }<<<3'd1 )+$signed( { 2'b0,x443 } <<<3'd1 )+$signed( { 2'b0,x699 } <<<3'd1 )-$signed(11'd16);
assign y45=temp_y[45][11] ==1'b1 ? 5'd0 :  
        temp_y[45][8] ==1'b1 ? 5'd31 : 
        temp_y[45][2]==1'b1 ? temp_y[45][7:3]+1'b1 : temp_y[45][7:3];
assign temp_y[109] = 
+$signed( { 3'b0,x170 }<<<3'd2 )+$signed( -{ 2'b0,x426 }<<<3'd1 )+$signed( -{ 2'b0,x682 }<<<3'd1 )+$signed( { 2'b0,x171 } <<<3'd1 )+$signed( -{ 3'b0,x427 }<<<3'd2)+$signed( { 1'b0,x683 }  )+$signed( -{ 1'b0,x186 } )+$signed( { 1'b0,x698 }  )+$signed( -{ 2'b0,x187 }<<<3'd1 )+$signed( -{ 1'b0,x443 } )+$signed( { 2'b0,x699 } <<<3'd1 )+$signed(11'd24);
assign y109=temp_y[109][11] ==1'b1 ? 5'd0 :  
        temp_y[109][8] ==1'b1 ? 5'd31 : 
        temp_y[109][2]==1'b1 ? temp_y[109][7:3]+1'b1 : temp_y[109][7:3];
assign temp_y[173] = 
+$signed( { 2'b0,x170 } <<<3'd1 )+$signed( { 2'b0,x426 } <<<3'd1 )+$signed( { 1'b0,x682 }  )+$signed( { 2'b0,x171 } <<<3'd1 )+$signed( -{ 1'b0,x427 } )+$signed( { 1'b0,x683 }  )+$signed( -{ 2'b0,x186 }<<<3'd1 )+$signed( -{ 2'b0,x442 }<<<3'd1 )+$signed( -{ 1'b0,x698 } )+$signed( -{ 1'b0,x187 } )+$signed( -{ 1'b0,x443 } )+$signed( -{ 1'b0,x699 } )+$signed(11'd16);
assign y173=temp_y[173][11] ==1'b1 ? 5'd0 :  
        temp_y[173][8] ==1'b1 ? 5'd31 : 
        temp_y[173][2]==1'b1 ? temp_y[173][7:3]+1'b1 : temp_y[173][7:3];
assign temp_y[237] = 
+$signed( { 1'b0,x170 }  )+$signed( -{ 1'b0,x426 } )+$signed( { 1'b0,x171 }  )+$signed( -{ 1'b0,x427 } )+$signed( { 2'b0,x186 } <<<3'd1 )+$signed( -{ 1'b0,x442 } )+$signed( -{ 1'b0,x698 } )+$signed( { 2'b0,x187 } <<<3'd1 )+$signed( -{ 1'b0,x443 } )+$signed( -{ 2'b0,x699 }<<<3'd1 )+$signed(11'd40);
assign y237=temp_y[237][11] ==1'b1 ? 5'd0 :  
        temp_y[237][8] ==1'b1 ? 5'd31 : 
        temp_y[237][2]==1'b1 ? temp_y[237][7:3]+1'b1 : temp_y[237][7:3];
assign temp_y[301] = 
+$signed( -{ 1'b0,x170 } )+$signed( { 2'b0,x426 } <<<3'd1 )+$signed( -{ 1'b0,x682 } )+$signed( -{ 1'b0,x171 } )+$signed( { 2'b0,x427 } <<<3'd1 )+$signed( -{ 2'b0,x683 }<<<3'd1 )+$signed( -{ 1'b0,x186 } )+$signed( { 2'b0,x442 } <<<3'd1 )+$signed( -{ 1'b0,x698 } )+$signed( -{ 2'b0,x187 }<<<3'd1 )+$signed( { 3'b0,x443 }<<<3'd2 )+$signed( -{ 2'b0,x699 }<<<3'd1 )+$signed(11'd32);
assign y301=temp_y[301][11] ==1'b1 ? 5'd0 :  
        temp_y[301][8] ==1'b1 ? 5'd31 : 
        temp_y[301][2]==1'b1 ? temp_y[301][7:3]+1'b1 : temp_y[301][7:3];
assign temp_y[365] = 
+$signed( -{ 1'b0,x170 } )+$signed( -{ 2'b0,x426 }<<<3'd1 )+$signed( -{ 1'b0,x682 } )+$signed( { 1'b0,x171 }  )+$signed( { 2'b0,x427 } <<<3'd1 )+$signed( { 1'b0,x683 }  )+$signed( { 1'b0,x186 }  )+$signed( { 2'b0,x442 } <<<3'd1 )+$signed( { 2'b0,x698 } <<<3'd1 )+$signed( -{ 1'b0,x187 } )+$signed( -{ 2'b0,x443 }<<<3'd1 )+$signed( -{ 1'b0,x699 } )-$signed(11'd68);
assign y365=temp_y[365][11] ==1'b1 ? 5'd0 :  
        temp_y[365][8] ==1'b1 ? 5'd31 : 
        temp_y[365][2]==1'b1 ? temp_y[365][7:3]+1'b1 : temp_y[365][7:3];
assign temp_y[429] = 
+$signed( { 1'b0,x426 }  )+$signed( { 1'b0,x683 }  )+$signed( { 1'b0,x699 }  )-$signed(11'd108);
assign y429=temp_y[429][11] ==1'b1 ? 5'd0 :  
        temp_y[429][8] ==1'b1 ? 5'd31 : 
        temp_y[429][2]==1'b1 ? temp_y[429][7:3]+1'b1 : temp_y[429][7:3];
assign temp_y[493] = 
+$signed( -{ 2'b0,x170 }<<<3'd1 )+$signed( { 2'b0,x682 } <<<3'd1 )+$signed( -{ 2'b0,x171 }<<<3'd1 )+$signed( { 1'b0,x427 }  )+$signed( { 1'b0,x683 }  )+$signed( -{ 2'b0,x186 }<<<3'd1 )+$signed( { 1'b0,x442 }  )+$signed( { 1'b0,x698 }  )+$signed( -{ 1'b0,x187 } )+$signed(11'd64);
assign y493=temp_y[493][11] ==1'b1 ? 5'd0 :  
        temp_y[493][8] ==1'b1 ? 5'd31 : 
        temp_y[493][2]==1'b1 ? temp_y[493][7:3]+1'b1 : temp_y[493][7:3];
assign temp_y[557] = 
+$signed( -{ 2'b0,x170 }<<<3'd1 )+$signed( -{ 1'b0,x426 } )+$signed( -{ 3'b0,x171 }<<<3'd2)+$signed( { 1'b0,x186 }  )+$signed( { 1'b0,x442 }  )+$signed( { 3'b0,x187 }<<<3'd2 )+$signed(11'd16);
assign y557=temp_y[557][11] ==1'b1 ? 5'd0 :  
        temp_y[557][8] ==1'b1 ? 5'd31 : 
        temp_y[557][2]==1'b1 ? temp_y[557][7:3]+1'b1 : temp_y[557][7:3];
assign temp_y[621] = 
+$signed( { 2'b0,x426 } <<<3'd1 )+$signed( { 2'b0,x682 } <<<3'd1 )+$signed( -{ 1'b0,x171 } )+$signed( -{ 2'b0,x427 }<<<3'd1 )+$signed( -{ 2'b0,x683 }<<<3'd1 )+$signed( { 2'b0,x442 } <<<3'd1 )+$signed( { 1'b0,x698 }  )+$signed( -{ 2'b0,x443 }<<<3'd1 )-$signed(11'd8);
assign y621=temp_y[621][11] ==1'b1 ? 5'd0 :  
        temp_y[621][8] ==1'b1 ? 5'd31 : 
        temp_y[621][2]==1'b1 ? temp_y[621][7:3]+1'b1 : temp_y[621][7:3];
assign temp_y[46] = 
+$signed( -{ 2'b0,x428 }<<<3'd1 )+$signed( -{ 1'b0,x684 } )+$signed( { 1'b0,x173 }  )+$signed( { 1'b0,x429 }  )+$signed( { 1'b0,x685 }  )+$signed( -{ 2'b0,x444 }<<<3'd1 )+$signed( -{ 2'b0,x700 }<<<3'd1 )+$signed( { 2'b0,x445 } <<<3'd1 )+$signed( { 2'b0,x701 } <<<3'd1 )-$signed(11'd16);
assign y46=temp_y[46][11] ==1'b1 ? 5'd0 :  
        temp_y[46][8] ==1'b1 ? 5'd31 : 
        temp_y[46][2]==1'b1 ? temp_y[46][7:3]+1'b1 : temp_y[46][7:3];
assign temp_y[110] = 
+$signed( { 3'b0,x172 }<<<3'd2 )+$signed( -{ 2'b0,x428 }<<<3'd1 )+$signed( -{ 2'b0,x684 }<<<3'd1 )+$signed( { 2'b0,x173 } <<<3'd1 )+$signed( -{ 3'b0,x429 }<<<3'd2)+$signed( { 1'b0,x685 }  )+$signed( -{ 1'b0,x188 } )+$signed( { 1'b0,x700 }  )+$signed( -{ 2'b0,x189 }<<<3'd1 )+$signed( -{ 1'b0,x445 } )+$signed( { 2'b0,x701 } <<<3'd1 )+$signed(11'd24);
assign y110=temp_y[110][11] ==1'b1 ? 5'd0 :  
        temp_y[110][8] ==1'b1 ? 5'd31 : 
        temp_y[110][2]==1'b1 ? temp_y[110][7:3]+1'b1 : temp_y[110][7:3];
assign temp_y[174] = 
+$signed( { 2'b0,x172 } <<<3'd1 )+$signed( { 2'b0,x428 } <<<3'd1 )+$signed( { 1'b0,x684 }  )+$signed( { 2'b0,x173 } <<<3'd1 )+$signed( -{ 1'b0,x429 } )+$signed( { 1'b0,x685 }  )+$signed( -{ 2'b0,x188 }<<<3'd1 )+$signed( -{ 2'b0,x444 }<<<3'd1 )+$signed( -{ 1'b0,x700 } )+$signed( -{ 1'b0,x189 } )+$signed( -{ 1'b0,x445 } )+$signed( -{ 1'b0,x701 } )+$signed(11'd16);
assign y174=temp_y[174][11] ==1'b1 ? 5'd0 :  
        temp_y[174][8] ==1'b1 ? 5'd31 : 
        temp_y[174][2]==1'b1 ? temp_y[174][7:3]+1'b1 : temp_y[174][7:3];
assign temp_y[238] = 
+$signed( { 1'b0,x172 }  )+$signed( -{ 1'b0,x428 } )+$signed( { 1'b0,x173 }  )+$signed( -{ 1'b0,x429 } )+$signed( { 2'b0,x188 } <<<3'd1 )+$signed( -{ 1'b0,x444 } )+$signed( -{ 1'b0,x700 } )+$signed( { 2'b0,x189 } <<<3'd1 )+$signed( -{ 1'b0,x445 } )+$signed( -{ 2'b0,x701 }<<<3'd1 )+$signed(11'd40);
assign y238=temp_y[238][11] ==1'b1 ? 5'd0 :  
        temp_y[238][8] ==1'b1 ? 5'd31 : 
        temp_y[238][2]==1'b1 ? temp_y[238][7:3]+1'b1 : temp_y[238][7:3];
assign temp_y[302] = 
+$signed( -{ 1'b0,x172 } )+$signed( { 2'b0,x428 } <<<3'd1 )+$signed( -{ 1'b0,x684 } )+$signed( -{ 1'b0,x173 } )+$signed( { 2'b0,x429 } <<<3'd1 )+$signed( -{ 2'b0,x685 }<<<3'd1 )+$signed( -{ 1'b0,x188 } )+$signed( { 2'b0,x444 } <<<3'd1 )+$signed( -{ 1'b0,x700 } )+$signed( -{ 2'b0,x189 }<<<3'd1 )+$signed( { 3'b0,x445 }<<<3'd2 )+$signed( -{ 2'b0,x701 }<<<3'd1 )+$signed(11'd32);
assign y302=temp_y[302][11] ==1'b1 ? 5'd0 :  
        temp_y[302][8] ==1'b1 ? 5'd31 : 
        temp_y[302][2]==1'b1 ? temp_y[302][7:3]+1'b1 : temp_y[302][7:3];
assign temp_y[366] = 
+$signed( -{ 1'b0,x172 } )+$signed( -{ 2'b0,x428 }<<<3'd1 )+$signed( -{ 1'b0,x684 } )+$signed( { 1'b0,x173 }  )+$signed( { 2'b0,x429 } <<<3'd1 )+$signed( { 1'b0,x685 }  )+$signed( { 1'b0,x188 }  )+$signed( { 2'b0,x444 } <<<3'd1 )+$signed( { 2'b0,x700 } <<<3'd1 )+$signed( -{ 1'b0,x189 } )+$signed( -{ 2'b0,x445 }<<<3'd1 )+$signed( -{ 1'b0,x701 } )-$signed(11'd68);
assign y366=temp_y[366][11] ==1'b1 ? 5'd0 :  
        temp_y[366][8] ==1'b1 ? 5'd31 : 
        temp_y[366][2]==1'b1 ? temp_y[366][7:3]+1'b1 : temp_y[366][7:3];
assign temp_y[430] = 
+$signed( { 1'b0,x428 }  )+$signed( { 1'b0,x685 }  )+$signed( { 1'b0,x701 }  )-$signed(11'd108);
assign y430=temp_y[430][11] ==1'b1 ? 5'd0 :  
        temp_y[430][8] ==1'b1 ? 5'd31 : 
        temp_y[430][2]==1'b1 ? temp_y[430][7:3]+1'b1 : temp_y[430][7:3];
assign temp_y[494] = 
+$signed( -{ 2'b0,x172 }<<<3'd1 )+$signed( { 2'b0,x684 } <<<3'd1 )+$signed( -{ 2'b0,x173 }<<<3'd1 )+$signed( { 1'b0,x429 }  )+$signed( { 1'b0,x685 }  )+$signed( -{ 2'b0,x188 }<<<3'd1 )+$signed( { 1'b0,x444 }  )+$signed( { 1'b0,x700 }  )+$signed( -{ 1'b0,x189 } )+$signed(11'd64);
assign y494=temp_y[494][11] ==1'b1 ? 5'd0 :  
        temp_y[494][8] ==1'b1 ? 5'd31 : 
        temp_y[494][2]==1'b1 ? temp_y[494][7:3]+1'b1 : temp_y[494][7:3];
assign temp_y[558] = 
+$signed( -{ 2'b0,x172 }<<<3'd1 )+$signed( -{ 1'b0,x428 } )+$signed( -{ 3'b0,x173 }<<<3'd2)+$signed( { 1'b0,x188 }  )+$signed( { 1'b0,x444 }  )+$signed( { 3'b0,x189 }<<<3'd2 )+$signed(11'd16);
assign y558=temp_y[558][11] ==1'b1 ? 5'd0 :  
        temp_y[558][8] ==1'b1 ? 5'd31 : 
        temp_y[558][2]==1'b1 ? temp_y[558][7:3]+1'b1 : temp_y[558][7:3];
assign temp_y[622] = 
+$signed( { 2'b0,x428 } <<<3'd1 )+$signed( { 2'b0,x684 } <<<3'd1 )+$signed( -{ 1'b0,x173 } )+$signed( -{ 2'b0,x429 }<<<3'd1 )+$signed( -{ 2'b0,x685 }<<<3'd1 )+$signed( { 2'b0,x444 } <<<3'd1 )+$signed( { 1'b0,x700 }  )+$signed( -{ 2'b0,x445 }<<<3'd1 )-$signed(11'd8);
assign y622=temp_y[622][11] ==1'b1 ? 5'd0 :  
        temp_y[622][8] ==1'b1 ? 5'd31 : 
        temp_y[622][2]==1'b1 ? temp_y[622][7:3]+1'b1 : temp_y[622][7:3];
assign temp_y[47] = 
+$signed( -{ 2'b0,x430 }<<<3'd1 )+$signed( -{ 1'b0,x686 } )+$signed( { 1'b0,x175 }  )+$signed( { 1'b0,x431 }  )+$signed( { 1'b0,x687 }  )+$signed( -{ 2'b0,x446 }<<<3'd1 )+$signed( -{ 2'b0,x702 }<<<3'd1 )+$signed( { 2'b0,x447 } <<<3'd1 )+$signed( { 2'b0,x703 } <<<3'd1 )-$signed(11'd16);
assign y47=temp_y[47][11] ==1'b1 ? 5'd0 :  
        temp_y[47][8] ==1'b1 ? 5'd31 : 
        temp_y[47][2]==1'b1 ? temp_y[47][7:3]+1'b1 : temp_y[47][7:3];
assign temp_y[111] = 
+$signed( { 3'b0,x174 }<<<3'd2 )+$signed( -{ 2'b0,x430 }<<<3'd1 )+$signed( -{ 2'b0,x686 }<<<3'd1 )+$signed( { 2'b0,x175 } <<<3'd1 )+$signed( -{ 3'b0,x431 }<<<3'd2)+$signed( { 1'b0,x687 }  )+$signed( -{ 1'b0,x190 } )+$signed( { 1'b0,x702 }  )+$signed( -{ 2'b0,x191 }<<<3'd1 )+$signed( -{ 1'b0,x447 } )+$signed( { 2'b0,x703 } <<<3'd1 )+$signed(11'd24);
assign y111=temp_y[111][11] ==1'b1 ? 5'd0 :  
        temp_y[111][8] ==1'b1 ? 5'd31 : 
        temp_y[111][2]==1'b1 ? temp_y[111][7:3]+1'b1 : temp_y[111][7:3];
assign temp_y[175] = 
+$signed( { 2'b0,x174 } <<<3'd1 )+$signed( { 2'b0,x430 } <<<3'd1 )+$signed( { 1'b0,x686 }  )+$signed( { 2'b0,x175 } <<<3'd1 )+$signed( -{ 1'b0,x431 } )+$signed( { 1'b0,x687 }  )+$signed( -{ 2'b0,x190 }<<<3'd1 )+$signed( -{ 2'b0,x446 }<<<3'd1 )+$signed( -{ 1'b0,x702 } )+$signed( -{ 1'b0,x191 } )+$signed( -{ 1'b0,x447 } )+$signed( -{ 1'b0,x703 } )+$signed(11'd16);
assign y175=temp_y[175][11] ==1'b1 ? 5'd0 :  
        temp_y[175][8] ==1'b1 ? 5'd31 : 
        temp_y[175][2]==1'b1 ? temp_y[175][7:3]+1'b1 : temp_y[175][7:3];
assign temp_y[239] = 
+$signed( { 1'b0,x174 }  )+$signed( -{ 1'b0,x430 } )+$signed( { 1'b0,x175 }  )+$signed( -{ 1'b0,x431 } )+$signed( { 2'b0,x190 } <<<3'd1 )+$signed( -{ 1'b0,x446 } )+$signed( -{ 1'b0,x702 } )+$signed( { 2'b0,x191 } <<<3'd1 )+$signed( -{ 1'b0,x447 } )+$signed( -{ 2'b0,x703 }<<<3'd1 )+$signed(11'd40);
assign y239=temp_y[239][11] ==1'b1 ? 5'd0 :  
        temp_y[239][8] ==1'b1 ? 5'd31 : 
        temp_y[239][2]==1'b1 ? temp_y[239][7:3]+1'b1 : temp_y[239][7:3];
assign temp_y[303] = 
+$signed( -{ 1'b0,x174 } )+$signed( { 2'b0,x430 } <<<3'd1 )+$signed( -{ 1'b0,x686 } )+$signed( -{ 1'b0,x175 } )+$signed( { 2'b0,x431 } <<<3'd1 )+$signed( -{ 2'b0,x687 }<<<3'd1 )+$signed( -{ 1'b0,x190 } )+$signed( { 2'b0,x446 } <<<3'd1 )+$signed( -{ 1'b0,x702 } )+$signed( -{ 2'b0,x191 }<<<3'd1 )+$signed( { 3'b0,x447 }<<<3'd2 )+$signed( -{ 2'b0,x703 }<<<3'd1 )+$signed(11'd32);
assign y303=temp_y[303][11] ==1'b1 ? 5'd0 :  
        temp_y[303][8] ==1'b1 ? 5'd31 : 
        temp_y[303][2]==1'b1 ? temp_y[303][7:3]+1'b1 : temp_y[303][7:3];
assign temp_y[367] = 
+$signed( -{ 1'b0,x174 } )+$signed( -{ 2'b0,x430 }<<<3'd1 )+$signed( -{ 1'b0,x686 } )+$signed( { 1'b0,x175 }  )+$signed( { 2'b0,x431 } <<<3'd1 )+$signed( { 1'b0,x687 }  )+$signed( { 1'b0,x190 }  )+$signed( { 2'b0,x446 } <<<3'd1 )+$signed( { 2'b0,x702 } <<<3'd1 )+$signed( -{ 1'b0,x191 } )+$signed( -{ 2'b0,x447 }<<<3'd1 )+$signed( -{ 1'b0,x703 } )-$signed(11'd68);
assign y367=temp_y[367][11] ==1'b1 ? 5'd0 :  
        temp_y[367][8] ==1'b1 ? 5'd31 : 
        temp_y[367][2]==1'b1 ? temp_y[367][7:3]+1'b1 : temp_y[367][7:3];
assign temp_y[431] = 
+$signed( { 1'b0,x430 }  )+$signed( { 1'b0,x687 }  )+$signed( { 1'b0,x703 }  )-$signed(11'd108);
assign y431=temp_y[431][11] ==1'b1 ? 5'd0 :  
        temp_y[431][8] ==1'b1 ? 5'd31 : 
        temp_y[431][2]==1'b1 ? temp_y[431][7:3]+1'b1 : temp_y[431][7:3];
assign temp_y[495] = 
+$signed( -{ 2'b0,x174 }<<<3'd1 )+$signed( { 2'b0,x686 } <<<3'd1 )+$signed( -{ 2'b0,x175 }<<<3'd1 )+$signed( { 1'b0,x431 }  )+$signed( { 1'b0,x687 }  )+$signed( -{ 2'b0,x190 }<<<3'd1 )+$signed( { 1'b0,x446 }  )+$signed( { 1'b0,x702 }  )+$signed( -{ 1'b0,x191 } )+$signed(11'd64);
assign y495=temp_y[495][11] ==1'b1 ? 5'd0 :  
        temp_y[495][8] ==1'b1 ? 5'd31 : 
        temp_y[495][2]==1'b1 ? temp_y[495][7:3]+1'b1 : temp_y[495][7:3];
assign temp_y[559] = 
+$signed( -{ 2'b0,x174 }<<<3'd1 )+$signed( -{ 1'b0,x430 } )+$signed( -{ 3'b0,x175 }<<<3'd2)+$signed( { 1'b0,x190 }  )+$signed( { 1'b0,x446 }  )+$signed( { 3'b0,x191 }<<<3'd2 )+$signed(11'd16);
assign y559=temp_y[559][11] ==1'b1 ? 5'd0 :  
        temp_y[559][8] ==1'b1 ? 5'd31 : 
        temp_y[559][2]==1'b1 ? temp_y[559][7:3]+1'b1 : temp_y[559][7:3];
assign temp_y[623] = 
+$signed( { 2'b0,x430 } <<<3'd1 )+$signed( { 2'b0,x686 } <<<3'd1 )+$signed( -{ 1'b0,x175 } )+$signed( -{ 2'b0,x431 }<<<3'd1 )+$signed( -{ 2'b0,x687 }<<<3'd1 )+$signed( { 2'b0,x446 } <<<3'd1 )+$signed( { 1'b0,x702 }  )+$signed( -{ 2'b0,x447 }<<<3'd1 )-$signed(11'd8);
assign y623=temp_y[623][11] ==1'b1 ? 5'd0 :  
        temp_y[623][8] ==1'b1 ? 5'd31 : 
        temp_y[623][2]==1'b1 ? temp_y[623][7:3]+1'b1 : temp_y[623][7:3];
assign temp_y[48] = 
+$signed( -{ 2'b0,x448 }<<<3'd1 )+$signed( -{ 1'b0,x704 } )+$signed( { 1'b0,x193 }  )+$signed( { 1'b0,x449 }  )+$signed( { 1'b0,x705 }  )+$signed( -{ 2'b0,x464 }<<<3'd1 )+$signed( -{ 2'b0,x720 }<<<3'd1 )+$signed( { 2'b0,x465 } <<<3'd1 )+$signed( { 2'b0,x721 } <<<3'd1 )-$signed(11'd16);
assign y48=temp_y[48][11] ==1'b1 ? 5'd0 :  
        temp_y[48][8] ==1'b1 ? 5'd31 : 
        temp_y[48][2]==1'b1 ? temp_y[48][7:3]+1'b1 : temp_y[48][7:3];
assign temp_y[112] = 
+$signed( { 3'b0,x192 }<<<3'd2 )+$signed( -{ 2'b0,x448 }<<<3'd1 )+$signed( -{ 2'b0,x704 }<<<3'd1 )+$signed( { 2'b0,x193 } <<<3'd1 )+$signed( -{ 3'b0,x449 }<<<3'd2)+$signed( { 1'b0,x705 }  )+$signed( -{ 1'b0,x208 } )+$signed( { 1'b0,x720 }  )+$signed( -{ 2'b0,x209 }<<<3'd1 )+$signed( -{ 1'b0,x465 } )+$signed( { 2'b0,x721 } <<<3'd1 )+$signed(11'd24);
assign y112=temp_y[112][11] ==1'b1 ? 5'd0 :  
        temp_y[112][8] ==1'b1 ? 5'd31 : 
        temp_y[112][2]==1'b1 ? temp_y[112][7:3]+1'b1 : temp_y[112][7:3];
assign temp_y[176] = 
+$signed( { 2'b0,x192 } <<<3'd1 )+$signed( { 2'b0,x448 } <<<3'd1 )+$signed( { 1'b0,x704 }  )+$signed( { 2'b0,x193 } <<<3'd1 )+$signed( -{ 1'b0,x449 } )+$signed( { 1'b0,x705 }  )+$signed( -{ 2'b0,x208 }<<<3'd1 )+$signed( -{ 2'b0,x464 }<<<3'd1 )+$signed( -{ 1'b0,x720 } )+$signed( -{ 1'b0,x209 } )+$signed( -{ 1'b0,x465 } )+$signed( -{ 1'b0,x721 } )+$signed(11'd16);
assign y176=temp_y[176][11] ==1'b1 ? 5'd0 :  
        temp_y[176][8] ==1'b1 ? 5'd31 : 
        temp_y[176][2]==1'b1 ? temp_y[176][7:3]+1'b1 : temp_y[176][7:3];
assign temp_y[240] = 
+$signed( { 1'b0,x192 }  )+$signed( -{ 1'b0,x448 } )+$signed( { 1'b0,x193 }  )+$signed( -{ 1'b0,x449 } )+$signed( { 2'b0,x208 } <<<3'd1 )+$signed( -{ 1'b0,x464 } )+$signed( -{ 1'b0,x720 } )+$signed( { 2'b0,x209 } <<<3'd1 )+$signed( -{ 1'b0,x465 } )+$signed( -{ 2'b0,x721 }<<<3'd1 )+$signed(11'd40);
assign y240=temp_y[240][11] ==1'b1 ? 5'd0 :  
        temp_y[240][8] ==1'b1 ? 5'd31 : 
        temp_y[240][2]==1'b1 ? temp_y[240][7:3]+1'b1 : temp_y[240][7:3];
assign temp_y[304] = 
+$signed( -{ 1'b0,x192 } )+$signed( { 2'b0,x448 } <<<3'd1 )+$signed( -{ 1'b0,x704 } )+$signed( -{ 1'b0,x193 } )+$signed( { 2'b0,x449 } <<<3'd1 )+$signed( -{ 2'b0,x705 }<<<3'd1 )+$signed( -{ 1'b0,x208 } )+$signed( { 2'b0,x464 } <<<3'd1 )+$signed( -{ 1'b0,x720 } )+$signed( -{ 2'b0,x209 }<<<3'd1 )+$signed( { 3'b0,x465 }<<<3'd2 )+$signed( -{ 2'b0,x721 }<<<3'd1 )+$signed(11'd32);
assign y304=temp_y[304][11] ==1'b1 ? 5'd0 :  
        temp_y[304][8] ==1'b1 ? 5'd31 : 
        temp_y[304][2]==1'b1 ? temp_y[304][7:3]+1'b1 : temp_y[304][7:3];
assign temp_y[368] = 
+$signed( -{ 1'b0,x192 } )+$signed( -{ 2'b0,x448 }<<<3'd1 )+$signed( -{ 1'b0,x704 } )+$signed( { 1'b0,x193 }  )+$signed( { 2'b0,x449 } <<<3'd1 )+$signed( { 1'b0,x705 }  )+$signed( { 1'b0,x208 }  )+$signed( { 2'b0,x464 } <<<3'd1 )+$signed( { 2'b0,x720 } <<<3'd1 )+$signed( -{ 1'b0,x209 } )+$signed( -{ 2'b0,x465 }<<<3'd1 )+$signed( -{ 1'b0,x721 } )-$signed(11'd68);
assign y368=temp_y[368][11] ==1'b1 ? 5'd0 :  
        temp_y[368][8] ==1'b1 ? 5'd31 : 
        temp_y[368][2]==1'b1 ? temp_y[368][7:3]+1'b1 : temp_y[368][7:3];
assign temp_y[432] = 
+$signed( { 1'b0,x448 }  )+$signed( { 1'b0,x705 }  )+$signed( { 1'b0,x721 }  )-$signed(11'd108);
assign y432=temp_y[432][11] ==1'b1 ? 5'd0 :  
        temp_y[432][8] ==1'b1 ? 5'd31 : 
        temp_y[432][2]==1'b1 ? temp_y[432][7:3]+1'b1 : temp_y[432][7:3];
assign temp_y[496] = 
+$signed( -{ 2'b0,x192 }<<<3'd1 )+$signed( { 2'b0,x704 } <<<3'd1 )+$signed( -{ 2'b0,x193 }<<<3'd1 )+$signed( { 1'b0,x449 }  )+$signed( { 1'b0,x705 }  )+$signed( -{ 2'b0,x208 }<<<3'd1 )+$signed( { 1'b0,x464 }  )+$signed( { 1'b0,x720 }  )+$signed( -{ 1'b0,x209 } )+$signed(11'd64);
assign y496=temp_y[496][11] ==1'b1 ? 5'd0 :  
        temp_y[496][8] ==1'b1 ? 5'd31 : 
        temp_y[496][2]==1'b1 ? temp_y[496][7:3]+1'b1 : temp_y[496][7:3];
assign temp_y[560] = 
+$signed( -{ 2'b0,x192 }<<<3'd1 )+$signed( -{ 1'b0,x448 } )+$signed( -{ 3'b0,x193 }<<<3'd2)+$signed( { 1'b0,x208 }  )+$signed( { 1'b0,x464 }  )+$signed( { 3'b0,x209 }<<<3'd2 )+$signed(11'd16);
assign y560=temp_y[560][11] ==1'b1 ? 5'd0 :  
        temp_y[560][8] ==1'b1 ? 5'd31 : 
        temp_y[560][2]==1'b1 ? temp_y[560][7:3]+1'b1 : temp_y[560][7:3];
assign temp_y[624] = 
+$signed( { 2'b0,x448 } <<<3'd1 )+$signed( { 2'b0,x704 } <<<3'd1 )+$signed( -{ 1'b0,x193 } )+$signed( -{ 2'b0,x449 }<<<3'd1 )+$signed( -{ 2'b0,x705 }<<<3'd1 )+$signed( { 2'b0,x464 } <<<3'd1 )+$signed( { 1'b0,x720 }  )+$signed( -{ 2'b0,x465 }<<<3'd1 )-$signed(11'd8);
assign y624=temp_y[624][11] ==1'b1 ? 5'd0 :  
        temp_y[624][8] ==1'b1 ? 5'd31 : 
        temp_y[624][2]==1'b1 ? temp_y[624][7:3]+1'b1 : temp_y[624][7:3];
assign temp_y[49] = 
+$signed( -{ 2'b0,x450 }<<<3'd1 )+$signed( -{ 1'b0,x706 } )+$signed( { 1'b0,x195 }  )+$signed( { 1'b0,x451 }  )+$signed( { 1'b0,x707 }  )+$signed( -{ 2'b0,x466 }<<<3'd1 )+$signed( -{ 2'b0,x722 }<<<3'd1 )+$signed( { 2'b0,x467 } <<<3'd1 )+$signed( { 2'b0,x723 } <<<3'd1 )-$signed(11'd16);
assign y49=temp_y[49][11] ==1'b1 ? 5'd0 :  
        temp_y[49][8] ==1'b1 ? 5'd31 : 
        temp_y[49][2]==1'b1 ? temp_y[49][7:3]+1'b1 : temp_y[49][7:3];
assign temp_y[113] = 
+$signed( { 3'b0,x194 }<<<3'd2 )+$signed( -{ 2'b0,x450 }<<<3'd1 )+$signed( -{ 2'b0,x706 }<<<3'd1 )+$signed( { 2'b0,x195 } <<<3'd1 )+$signed( -{ 3'b0,x451 }<<<3'd2)+$signed( { 1'b0,x707 }  )+$signed( -{ 1'b0,x210 } )+$signed( { 1'b0,x722 }  )+$signed( -{ 2'b0,x211 }<<<3'd1 )+$signed( -{ 1'b0,x467 } )+$signed( { 2'b0,x723 } <<<3'd1 )+$signed(11'd24);
assign y113=temp_y[113][11] ==1'b1 ? 5'd0 :  
        temp_y[113][8] ==1'b1 ? 5'd31 : 
        temp_y[113][2]==1'b1 ? temp_y[113][7:3]+1'b1 : temp_y[113][7:3];
assign temp_y[177] = 
+$signed( { 2'b0,x194 } <<<3'd1 )+$signed( { 2'b0,x450 } <<<3'd1 )+$signed( { 1'b0,x706 }  )+$signed( { 2'b0,x195 } <<<3'd1 )+$signed( -{ 1'b0,x451 } )+$signed( { 1'b0,x707 }  )+$signed( -{ 2'b0,x210 }<<<3'd1 )+$signed( -{ 2'b0,x466 }<<<3'd1 )+$signed( -{ 1'b0,x722 } )+$signed( -{ 1'b0,x211 } )+$signed( -{ 1'b0,x467 } )+$signed( -{ 1'b0,x723 } )+$signed(11'd16);
assign y177=temp_y[177][11] ==1'b1 ? 5'd0 :  
        temp_y[177][8] ==1'b1 ? 5'd31 : 
        temp_y[177][2]==1'b1 ? temp_y[177][7:3]+1'b1 : temp_y[177][7:3];
assign temp_y[241] = 
+$signed( { 1'b0,x194 }  )+$signed( -{ 1'b0,x450 } )+$signed( { 1'b0,x195 }  )+$signed( -{ 1'b0,x451 } )+$signed( { 2'b0,x210 } <<<3'd1 )+$signed( -{ 1'b0,x466 } )+$signed( -{ 1'b0,x722 } )+$signed( { 2'b0,x211 } <<<3'd1 )+$signed( -{ 1'b0,x467 } )+$signed( -{ 2'b0,x723 }<<<3'd1 )+$signed(11'd40);
assign y241=temp_y[241][11] ==1'b1 ? 5'd0 :  
        temp_y[241][8] ==1'b1 ? 5'd31 : 
        temp_y[241][2]==1'b1 ? temp_y[241][7:3]+1'b1 : temp_y[241][7:3];
assign temp_y[305] = 
+$signed( -{ 1'b0,x194 } )+$signed( { 2'b0,x450 } <<<3'd1 )+$signed( -{ 1'b0,x706 } )+$signed( -{ 1'b0,x195 } )+$signed( { 2'b0,x451 } <<<3'd1 )+$signed( -{ 2'b0,x707 }<<<3'd1 )+$signed( -{ 1'b0,x210 } )+$signed( { 2'b0,x466 } <<<3'd1 )+$signed( -{ 1'b0,x722 } )+$signed( -{ 2'b0,x211 }<<<3'd1 )+$signed( { 3'b0,x467 }<<<3'd2 )+$signed( -{ 2'b0,x723 }<<<3'd1 )+$signed(11'd32);
assign y305=temp_y[305][11] ==1'b1 ? 5'd0 :  
        temp_y[305][8] ==1'b1 ? 5'd31 : 
        temp_y[305][2]==1'b1 ? temp_y[305][7:3]+1'b1 : temp_y[305][7:3];
assign temp_y[369] = 
+$signed( -{ 1'b0,x194 } )+$signed( -{ 2'b0,x450 }<<<3'd1 )+$signed( -{ 1'b0,x706 } )+$signed( { 1'b0,x195 }  )+$signed( { 2'b0,x451 } <<<3'd1 )+$signed( { 1'b0,x707 }  )+$signed( { 1'b0,x210 }  )+$signed( { 2'b0,x466 } <<<3'd1 )+$signed( { 2'b0,x722 } <<<3'd1 )+$signed( -{ 1'b0,x211 } )+$signed( -{ 2'b0,x467 }<<<3'd1 )+$signed( -{ 1'b0,x723 } )-$signed(11'd68);
assign y369=temp_y[369][11] ==1'b1 ? 5'd0 :  
        temp_y[369][8] ==1'b1 ? 5'd31 : 
        temp_y[369][2]==1'b1 ? temp_y[369][7:3]+1'b1 : temp_y[369][7:3];
assign temp_y[433] = 
+$signed( { 1'b0,x450 }  )+$signed( { 1'b0,x707 }  )+$signed( { 1'b0,x723 }  )-$signed(11'd108);
assign y433=temp_y[433][11] ==1'b1 ? 5'd0 :  
        temp_y[433][8] ==1'b1 ? 5'd31 : 
        temp_y[433][2]==1'b1 ? temp_y[433][7:3]+1'b1 : temp_y[433][7:3];
assign temp_y[497] = 
+$signed( -{ 2'b0,x194 }<<<3'd1 )+$signed( { 2'b0,x706 } <<<3'd1 )+$signed( -{ 2'b0,x195 }<<<3'd1 )+$signed( { 1'b0,x451 }  )+$signed( { 1'b0,x707 }  )+$signed( -{ 2'b0,x210 }<<<3'd1 )+$signed( { 1'b0,x466 }  )+$signed( { 1'b0,x722 }  )+$signed( -{ 1'b0,x211 } )+$signed(11'd64);
assign y497=temp_y[497][11] ==1'b1 ? 5'd0 :  
        temp_y[497][8] ==1'b1 ? 5'd31 : 
        temp_y[497][2]==1'b1 ? temp_y[497][7:3]+1'b1 : temp_y[497][7:3];
assign temp_y[561] = 
+$signed( -{ 2'b0,x194 }<<<3'd1 )+$signed( -{ 1'b0,x450 } )+$signed( -{ 3'b0,x195 }<<<3'd2)+$signed( { 1'b0,x210 }  )+$signed( { 1'b0,x466 }  )+$signed( { 3'b0,x211 }<<<3'd2 )+$signed(11'd16);
assign y561=temp_y[561][11] ==1'b1 ? 5'd0 :  
        temp_y[561][8] ==1'b1 ? 5'd31 : 
        temp_y[561][2]==1'b1 ? temp_y[561][7:3]+1'b1 : temp_y[561][7:3];
assign temp_y[625] = 
+$signed( { 2'b0,x450 } <<<3'd1 )+$signed( { 2'b0,x706 } <<<3'd1 )+$signed( -{ 1'b0,x195 } )+$signed( -{ 2'b0,x451 }<<<3'd1 )+$signed( -{ 2'b0,x707 }<<<3'd1 )+$signed( { 2'b0,x466 } <<<3'd1 )+$signed( { 1'b0,x722 }  )+$signed( -{ 2'b0,x467 }<<<3'd1 )-$signed(11'd8);
assign y625=temp_y[625][11] ==1'b1 ? 5'd0 :  
        temp_y[625][8] ==1'b1 ? 5'd31 : 
        temp_y[625][2]==1'b1 ? temp_y[625][7:3]+1'b1 : temp_y[625][7:3];
assign temp_y[50] = 
+$signed( -{ 2'b0,x452 }<<<3'd1 )+$signed( -{ 1'b0,x708 } )+$signed( { 1'b0,x197 }  )+$signed( { 1'b0,x453 }  )+$signed( { 1'b0,x709 }  )+$signed( -{ 2'b0,x468 }<<<3'd1 )+$signed( -{ 2'b0,x724 }<<<3'd1 )+$signed( { 2'b0,x469 } <<<3'd1 )+$signed( { 2'b0,x725 } <<<3'd1 )-$signed(11'd16);
assign y50=temp_y[50][11] ==1'b1 ? 5'd0 :  
        temp_y[50][8] ==1'b1 ? 5'd31 : 
        temp_y[50][2]==1'b1 ? temp_y[50][7:3]+1'b1 : temp_y[50][7:3];
assign temp_y[114] = 
+$signed( { 3'b0,x196 }<<<3'd2 )+$signed( -{ 2'b0,x452 }<<<3'd1 )+$signed( -{ 2'b0,x708 }<<<3'd1 )+$signed( { 2'b0,x197 } <<<3'd1 )+$signed( -{ 3'b0,x453 }<<<3'd2)+$signed( { 1'b0,x709 }  )+$signed( -{ 1'b0,x212 } )+$signed( { 1'b0,x724 }  )+$signed( -{ 2'b0,x213 }<<<3'd1 )+$signed( -{ 1'b0,x469 } )+$signed( { 2'b0,x725 } <<<3'd1 )+$signed(11'd24);
assign y114=temp_y[114][11] ==1'b1 ? 5'd0 :  
        temp_y[114][8] ==1'b1 ? 5'd31 : 
        temp_y[114][2]==1'b1 ? temp_y[114][7:3]+1'b1 : temp_y[114][7:3];
assign temp_y[178] = 
+$signed( { 2'b0,x196 } <<<3'd1 )+$signed( { 2'b0,x452 } <<<3'd1 )+$signed( { 1'b0,x708 }  )+$signed( { 2'b0,x197 } <<<3'd1 )+$signed( -{ 1'b0,x453 } )+$signed( { 1'b0,x709 }  )+$signed( -{ 2'b0,x212 }<<<3'd1 )+$signed( -{ 2'b0,x468 }<<<3'd1 )+$signed( -{ 1'b0,x724 } )+$signed( -{ 1'b0,x213 } )+$signed( -{ 1'b0,x469 } )+$signed( -{ 1'b0,x725 } )+$signed(11'd16);
assign y178=temp_y[178][11] ==1'b1 ? 5'd0 :  
        temp_y[178][8] ==1'b1 ? 5'd31 : 
        temp_y[178][2]==1'b1 ? temp_y[178][7:3]+1'b1 : temp_y[178][7:3];
assign temp_y[242] = 
+$signed( { 1'b0,x196 }  )+$signed( -{ 1'b0,x452 } )+$signed( { 1'b0,x197 }  )+$signed( -{ 1'b0,x453 } )+$signed( { 2'b0,x212 } <<<3'd1 )+$signed( -{ 1'b0,x468 } )+$signed( -{ 1'b0,x724 } )+$signed( { 2'b0,x213 } <<<3'd1 )+$signed( -{ 1'b0,x469 } )+$signed( -{ 2'b0,x725 }<<<3'd1 )+$signed(11'd40);
assign y242=temp_y[242][11] ==1'b1 ? 5'd0 :  
        temp_y[242][8] ==1'b1 ? 5'd31 : 
        temp_y[242][2]==1'b1 ? temp_y[242][7:3]+1'b1 : temp_y[242][7:3];
assign temp_y[306] = 
+$signed( -{ 1'b0,x196 } )+$signed( { 2'b0,x452 } <<<3'd1 )+$signed( -{ 1'b0,x708 } )+$signed( -{ 1'b0,x197 } )+$signed( { 2'b0,x453 } <<<3'd1 )+$signed( -{ 2'b0,x709 }<<<3'd1 )+$signed( -{ 1'b0,x212 } )+$signed( { 2'b0,x468 } <<<3'd1 )+$signed( -{ 1'b0,x724 } )+$signed( -{ 2'b0,x213 }<<<3'd1 )+$signed( { 3'b0,x469 }<<<3'd2 )+$signed( -{ 2'b0,x725 }<<<3'd1 )+$signed(11'd32);
assign y306=temp_y[306][11] ==1'b1 ? 5'd0 :  
        temp_y[306][8] ==1'b1 ? 5'd31 : 
        temp_y[306][2]==1'b1 ? temp_y[306][7:3]+1'b1 : temp_y[306][7:3];
assign temp_y[370] = 
+$signed( -{ 1'b0,x196 } )+$signed( -{ 2'b0,x452 }<<<3'd1 )+$signed( -{ 1'b0,x708 } )+$signed( { 1'b0,x197 }  )+$signed( { 2'b0,x453 } <<<3'd1 )+$signed( { 1'b0,x709 }  )+$signed( { 1'b0,x212 }  )+$signed( { 2'b0,x468 } <<<3'd1 )+$signed( { 2'b0,x724 } <<<3'd1 )+$signed( -{ 1'b0,x213 } )+$signed( -{ 2'b0,x469 }<<<3'd1 )+$signed( -{ 1'b0,x725 } )-$signed(11'd68);
assign y370=temp_y[370][11] ==1'b1 ? 5'd0 :  
        temp_y[370][8] ==1'b1 ? 5'd31 : 
        temp_y[370][2]==1'b1 ? temp_y[370][7:3]+1'b1 : temp_y[370][7:3];
assign temp_y[434] = 
+$signed( { 1'b0,x452 }  )+$signed( { 1'b0,x709 }  )+$signed( { 1'b0,x725 }  )-$signed(11'd108);
assign y434=temp_y[434][11] ==1'b1 ? 5'd0 :  
        temp_y[434][8] ==1'b1 ? 5'd31 : 
        temp_y[434][2]==1'b1 ? temp_y[434][7:3]+1'b1 : temp_y[434][7:3];
assign temp_y[498] = 
+$signed( -{ 2'b0,x196 }<<<3'd1 )+$signed( { 2'b0,x708 } <<<3'd1 )+$signed( -{ 2'b0,x197 }<<<3'd1 )+$signed( { 1'b0,x453 }  )+$signed( { 1'b0,x709 }  )+$signed( -{ 2'b0,x212 }<<<3'd1 )+$signed( { 1'b0,x468 }  )+$signed( { 1'b0,x724 }  )+$signed( -{ 1'b0,x213 } )+$signed(11'd64);
assign y498=temp_y[498][11] ==1'b1 ? 5'd0 :  
        temp_y[498][8] ==1'b1 ? 5'd31 : 
        temp_y[498][2]==1'b1 ? temp_y[498][7:3]+1'b1 : temp_y[498][7:3];
assign temp_y[562] = 
+$signed( -{ 2'b0,x196 }<<<3'd1 )+$signed( -{ 1'b0,x452 } )+$signed( -{ 3'b0,x197 }<<<3'd2)+$signed( { 1'b0,x212 }  )+$signed( { 1'b0,x468 }  )+$signed( { 3'b0,x213 }<<<3'd2 )+$signed(11'd16);
assign y562=temp_y[562][11] ==1'b1 ? 5'd0 :  
        temp_y[562][8] ==1'b1 ? 5'd31 : 
        temp_y[562][2]==1'b1 ? temp_y[562][7:3]+1'b1 : temp_y[562][7:3];
assign temp_y[626] = 
+$signed( { 2'b0,x452 } <<<3'd1 )+$signed( { 2'b0,x708 } <<<3'd1 )+$signed( -{ 1'b0,x197 } )+$signed( -{ 2'b0,x453 }<<<3'd1 )+$signed( -{ 2'b0,x709 }<<<3'd1 )+$signed( { 2'b0,x468 } <<<3'd1 )+$signed( { 1'b0,x724 }  )+$signed( -{ 2'b0,x469 }<<<3'd1 )-$signed(11'd8);
assign y626=temp_y[626][11] ==1'b1 ? 5'd0 :  
        temp_y[626][8] ==1'b1 ? 5'd31 : 
        temp_y[626][2]==1'b1 ? temp_y[626][7:3]+1'b1 : temp_y[626][7:3];
assign temp_y[51] = 
+$signed( -{ 2'b0,x454 }<<<3'd1 )+$signed( -{ 1'b0,x710 } )+$signed( { 1'b0,x199 }  )+$signed( { 1'b0,x455 }  )+$signed( { 1'b0,x711 }  )+$signed( -{ 2'b0,x470 }<<<3'd1 )+$signed( -{ 2'b0,x726 }<<<3'd1 )+$signed( { 2'b0,x471 } <<<3'd1 )+$signed( { 2'b0,x727 } <<<3'd1 )-$signed(11'd16);
assign y51=temp_y[51][11] ==1'b1 ? 5'd0 :  
        temp_y[51][8] ==1'b1 ? 5'd31 : 
        temp_y[51][2]==1'b1 ? temp_y[51][7:3]+1'b1 : temp_y[51][7:3];
assign temp_y[115] = 
+$signed( { 3'b0,x198 }<<<3'd2 )+$signed( -{ 2'b0,x454 }<<<3'd1 )+$signed( -{ 2'b0,x710 }<<<3'd1 )+$signed( { 2'b0,x199 } <<<3'd1 )+$signed( -{ 3'b0,x455 }<<<3'd2)+$signed( { 1'b0,x711 }  )+$signed( -{ 1'b0,x214 } )+$signed( { 1'b0,x726 }  )+$signed( -{ 2'b0,x215 }<<<3'd1 )+$signed( -{ 1'b0,x471 } )+$signed( { 2'b0,x727 } <<<3'd1 )+$signed(11'd24);
assign y115=temp_y[115][11] ==1'b1 ? 5'd0 :  
        temp_y[115][8] ==1'b1 ? 5'd31 : 
        temp_y[115][2]==1'b1 ? temp_y[115][7:3]+1'b1 : temp_y[115][7:3];
assign temp_y[179] = 
+$signed( { 2'b0,x198 } <<<3'd1 )+$signed( { 2'b0,x454 } <<<3'd1 )+$signed( { 1'b0,x710 }  )+$signed( { 2'b0,x199 } <<<3'd1 )+$signed( -{ 1'b0,x455 } )+$signed( { 1'b0,x711 }  )+$signed( -{ 2'b0,x214 }<<<3'd1 )+$signed( -{ 2'b0,x470 }<<<3'd1 )+$signed( -{ 1'b0,x726 } )+$signed( -{ 1'b0,x215 } )+$signed( -{ 1'b0,x471 } )+$signed( -{ 1'b0,x727 } )+$signed(11'd16);
assign y179=temp_y[179][11] ==1'b1 ? 5'd0 :  
        temp_y[179][8] ==1'b1 ? 5'd31 : 
        temp_y[179][2]==1'b1 ? temp_y[179][7:3]+1'b1 : temp_y[179][7:3];
assign temp_y[243] = 
+$signed( { 1'b0,x198 }  )+$signed( -{ 1'b0,x454 } )+$signed( { 1'b0,x199 }  )+$signed( -{ 1'b0,x455 } )+$signed( { 2'b0,x214 } <<<3'd1 )+$signed( -{ 1'b0,x470 } )+$signed( -{ 1'b0,x726 } )+$signed( { 2'b0,x215 } <<<3'd1 )+$signed( -{ 1'b0,x471 } )+$signed( -{ 2'b0,x727 }<<<3'd1 )+$signed(11'd40);
assign y243=temp_y[243][11] ==1'b1 ? 5'd0 :  
        temp_y[243][8] ==1'b1 ? 5'd31 : 
        temp_y[243][2]==1'b1 ? temp_y[243][7:3]+1'b1 : temp_y[243][7:3];
assign temp_y[307] = 
+$signed( -{ 1'b0,x198 } )+$signed( { 2'b0,x454 } <<<3'd1 )+$signed( -{ 1'b0,x710 } )+$signed( -{ 1'b0,x199 } )+$signed( { 2'b0,x455 } <<<3'd1 )+$signed( -{ 2'b0,x711 }<<<3'd1 )+$signed( -{ 1'b0,x214 } )+$signed( { 2'b0,x470 } <<<3'd1 )+$signed( -{ 1'b0,x726 } )+$signed( -{ 2'b0,x215 }<<<3'd1 )+$signed( { 3'b0,x471 }<<<3'd2 )+$signed( -{ 2'b0,x727 }<<<3'd1 )+$signed(11'd32);
assign y307=temp_y[307][11] ==1'b1 ? 5'd0 :  
        temp_y[307][8] ==1'b1 ? 5'd31 : 
        temp_y[307][2]==1'b1 ? temp_y[307][7:3]+1'b1 : temp_y[307][7:3];
assign temp_y[371] = 
+$signed( -{ 1'b0,x198 } )+$signed( -{ 2'b0,x454 }<<<3'd1 )+$signed( -{ 1'b0,x710 } )+$signed( { 1'b0,x199 }  )+$signed( { 2'b0,x455 } <<<3'd1 )+$signed( { 1'b0,x711 }  )+$signed( { 1'b0,x214 }  )+$signed( { 2'b0,x470 } <<<3'd1 )+$signed( { 2'b0,x726 } <<<3'd1 )+$signed( -{ 1'b0,x215 } )+$signed( -{ 2'b0,x471 }<<<3'd1 )+$signed( -{ 1'b0,x727 } )-$signed(11'd68);
assign y371=temp_y[371][11] ==1'b1 ? 5'd0 :  
        temp_y[371][8] ==1'b1 ? 5'd31 : 
        temp_y[371][2]==1'b1 ? temp_y[371][7:3]+1'b1 : temp_y[371][7:3];
assign temp_y[435] = 
+$signed( { 1'b0,x454 }  )+$signed( { 1'b0,x711 }  )+$signed( { 1'b0,x727 }  )-$signed(11'd108);
assign y435=temp_y[435][11] ==1'b1 ? 5'd0 :  
        temp_y[435][8] ==1'b1 ? 5'd31 : 
        temp_y[435][2]==1'b1 ? temp_y[435][7:3]+1'b1 : temp_y[435][7:3];
assign temp_y[499] = 
+$signed( -{ 2'b0,x198 }<<<3'd1 )+$signed( { 2'b0,x710 } <<<3'd1 )+$signed( -{ 2'b0,x199 }<<<3'd1 )+$signed( { 1'b0,x455 }  )+$signed( { 1'b0,x711 }  )+$signed( -{ 2'b0,x214 }<<<3'd1 )+$signed( { 1'b0,x470 }  )+$signed( { 1'b0,x726 }  )+$signed( -{ 1'b0,x215 } )+$signed(11'd64);
assign y499=temp_y[499][11] ==1'b1 ? 5'd0 :  
        temp_y[499][8] ==1'b1 ? 5'd31 : 
        temp_y[499][2]==1'b1 ? temp_y[499][7:3]+1'b1 : temp_y[499][7:3];
assign temp_y[563] = 
+$signed( -{ 2'b0,x198 }<<<3'd1 )+$signed( -{ 1'b0,x454 } )+$signed( -{ 3'b0,x199 }<<<3'd2)+$signed( { 1'b0,x214 }  )+$signed( { 1'b0,x470 }  )+$signed( { 3'b0,x215 }<<<3'd2 )+$signed(11'd16);
assign y563=temp_y[563][11] ==1'b1 ? 5'd0 :  
        temp_y[563][8] ==1'b1 ? 5'd31 : 
        temp_y[563][2]==1'b1 ? temp_y[563][7:3]+1'b1 : temp_y[563][7:3];
assign temp_y[627] = 
+$signed( { 2'b0,x454 } <<<3'd1 )+$signed( { 2'b0,x710 } <<<3'd1 )+$signed( -{ 1'b0,x199 } )+$signed( -{ 2'b0,x455 }<<<3'd1 )+$signed( -{ 2'b0,x711 }<<<3'd1 )+$signed( { 2'b0,x470 } <<<3'd1 )+$signed( { 1'b0,x726 }  )+$signed( -{ 2'b0,x471 }<<<3'd1 )-$signed(11'd8);
assign y627=temp_y[627][11] ==1'b1 ? 5'd0 :  
        temp_y[627][8] ==1'b1 ? 5'd31 : 
        temp_y[627][2]==1'b1 ? temp_y[627][7:3]+1'b1 : temp_y[627][7:3];
assign temp_y[52] = 
+$signed( -{ 2'b0,x456 }<<<3'd1 )+$signed( -{ 1'b0,x712 } )+$signed( { 1'b0,x201 }  )+$signed( { 1'b0,x457 }  )+$signed( { 1'b0,x713 }  )+$signed( -{ 2'b0,x472 }<<<3'd1 )+$signed( -{ 2'b0,x728 }<<<3'd1 )+$signed( { 2'b0,x473 } <<<3'd1 )+$signed( { 2'b0,x729 } <<<3'd1 )-$signed(11'd16);
assign y52=temp_y[52][11] ==1'b1 ? 5'd0 :  
        temp_y[52][8] ==1'b1 ? 5'd31 : 
        temp_y[52][2]==1'b1 ? temp_y[52][7:3]+1'b1 : temp_y[52][7:3];
assign temp_y[116] = 
+$signed( { 3'b0,x200 }<<<3'd2 )+$signed( -{ 2'b0,x456 }<<<3'd1 )+$signed( -{ 2'b0,x712 }<<<3'd1 )+$signed( { 2'b0,x201 } <<<3'd1 )+$signed( -{ 3'b0,x457 }<<<3'd2)+$signed( { 1'b0,x713 }  )+$signed( -{ 1'b0,x216 } )+$signed( { 1'b0,x728 }  )+$signed( -{ 2'b0,x217 }<<<3'd1 )+$signed( -{ 1'b0,x473 } )+$signed( { 2'b0,x729 } <<<3'd1 )+$signed(11'd24);
assign y116=temp_y[116][11] ==1'b1 ? 5'd0 :  
        temp_y[116][8] ==1'b1 ? 5'd31 : 
        temp_y[116][2]==1'b1 ? temp_y[116][7:3]+1'b1 : temp_y[116][7:3];
assign temp_y[180] = 
+$signed( { 2'b0,x200 } <<<3'd1 )+$signed( { 2'b0,x456 } <<<3'd1 )+$signed( { 1'b0,x712 }  )+$signed( { 2'b0,x201 } <<<3'd1 )+$signed( -{ 1'b0,x457 } )+$signed( { 1'b0,x713 }  )+$signed( -{ 2'b0,x216 }<<<3'd1 )+$signed( -{ 2'b0,x472 }<<<3'd1 )+$signed( -{ 1'b0,x728 } )+$signed( -{ 1'b0,x217 } )+$signed( -{ 1'b0,x473 } )+$signed( -{ 1'b0,x729 } )+$signed(11'd16);
assign y180=temp_y[180][11] ==1'b1 ? 5'd0 :  
        temp_y[180][8] ==1'b1 ? 5'd31 : 
        temp_y[180][2]==1'b1 ? temp_y[180][7:3]+1'b1 : temp_y[180][7:3];
assign temp_y[244] = 
+$signed( { 1'b0,x200 }  )+$signed( -{ 1'b0,x456 } )+$signed( { 1'b0,x201 }  )+$signed( -{ 1'b0,x457 } )+$signed( { 2'b0,x216 } <<<3'd1 )+$signed( -{ 1'b0,x472 } )+$signed( -{ 1'b0,x728 } )+$signed( { 2'b0,x217 } <<<3'd1 )+$signed( -{ 1'b0,x473 } )+$signed( -{ 2'b0,x729 }<<<3'd1 )+$signed(11'd40);
assign y244=temp_y[244][11] ==1'b1 ? 5'd0 :  
        temp_y[244][8] ==1'b1 ? 5'd31 : 
        temp_y[244][2]==1'b1 ? temp_y[244][7:3]+1'b1 : temp_y[244][7:3];
assign temp_y[308] = 
+$signed( -{ 1'b0,x200 } )+$signed( { 2'b0,x456 } <<<3'd1 )+$signed( -{ 1'b0,x712 } )+$signed( -{ 1'b0,x201 } )+$signed( { 2'b0,x457 } <<<3'd1 )+$signed( -{ 2'b0,x713 }<<<3'd1 )+$signed( -{ 1'b0,x216 } )+$signed( { 2'b0,x472 } <<<3'd1 )+$signed( -{ 1'b0,x728 } )+$signed( -{ 2'b0,x217 }<<<3'd1 )+$signed( { 3'b0,x473 }<<<3'd2 )+$signed( -{ 2'b0,x729 }<<<3'd1 )+$signed(11'd32);
assign y308=temp_y[308][11] ==1'b1 ? 5'd0 :  
        temp_y[308][8] ==1'b1 ? 5'd31 : 
        temp_y[308][2]==1'b1 ? temp_y[308][7:3]+1'b1 : temp_y[308][7:3];
assign temp_y[372] = 
+$signed( -{ 1'b0,x200 } )+$signed( -{ 2'b0,x456 }<<<3'd1 )+$signed( -{ 1'b0,x712 } )+$signed( { 1'b0,x201 }  )+$signed( { 2'b0,x457 } <<<3'd1 )+$signed( { 1'b0,x713 }  )+$signed( { 1'b0,x216 }  )+$signed( { 2'b0,x472 } <<<3'd1 )+$signed( { 2'b0,x728 } <<<3'd1 )+$signed( -{ 1'b0,x217 } )+$signed( -{ 2'b0,x473 }<<<3'd1 )+$signed( -{ 1'b0,x729 } )-$signed(11'd68);
assign y372=temp_y[372][11] ==1'b1 ? 5'd0 :  
        temp_y[372][8] ==1'b1 ? 5'd31 : 
        temp_y[372][2]==1'b1 ? temp_y[372][7:3]+1'b1 : temp_y[372][7:3];
assign temp_y[436] = 
+$signed( { 1'b0,x456 }  )+$signed( { 1'b0,x713 }  )+$signed( { 1'b0,x729 }  )-$signed(11'd108);
assign y436=temp_y[436][11] ==1'b1 ? 5'd0 :  
        temp_y[436][8] ==1'b1 ? 5'd31 : 
        temp_y[436][2]==1'b1 ? temp_y[436][7:3]+1'b1 : temp_y[436][7:3];
assign temp_y[500] = 
+$signed( -{ 2'b0,x200 }<<<3'd1 )+$signed( { 2'b0,x712 } <<<3'd1 )+$signed( -{ 2'b0,x201 }<<<3'd1 )+$signed( { 1'b0,x457 }  )+$signed( { 1'b0,x713 }  )+$signed( -{ 2'b0,x216 }<<<3'd1 )+$signed( { 1'b0,x472 }  )+$signed( { 1'b0,x728 }  )+$signed( -{ 1'b0,x217 } )+$signed(11'd64);
assign y500=temp_y[500][11] ==1'b1 ? 5'd0 :  
        temp_y[500][8] ==1'b1 ? 5'd31 : 
        temp_y[500][2]==1'b1 ? temp_y[500][7:3]+1'b1 : temp_y[500][7:3];
assign temp_y[564] = 
+$signed( -{ 2'b0,x200 }<<<3'd1 )+$signed( -{ 1'b0,x456 } )+$signed( -{ 3'b0,x201 }<<<3'd2)+$signed( { 1'b0,x216 }  )+$signed( { 1'b0,x472 }  )+$signed( { 3'b0,x217 }<<<3'd2 )+$signed(11'd16);
assign y564=temp_y[564][11] ==1'b1 ? 5'd0 :  
        temp_y[564][8] ==1'b1 ? 5'd31 : 
        temp_y[564][2]==1'b1 ? temp_y[564][7:3]+1'b1 : temp_y[564][7:3];
assign temp_y[628] = 
+$signed( { 2'b0,x456 } <<<3'd1 )+$signed( { 2'b0,x712 } <<<3'd1 )+$signed( -{ 1'b0,x201 } )+$signed( -{ 2'b0,x457 }<<<3'd1 )+$signed( -{ 2'b0,x713 }<<<3'd1 )+$signed( { 2'b0,x472 } <<<3'd1 )+$signed( { 1'b0,x728 }  )+$signed( -{ 2'b0,x473 }<<<3'd1 )-$signed(11'd8);
assign y628=temp_y[628][11] ==1'b1 ? 5'd0 :  
        temp_y[628][8] ==1'b1 ? 5'd31 : 
        temp_y[628][2]==1'b1 ? temp_y[628][7:3]+1'b1 : temp_y[628][7:3];
assign temp_y[53] = 
+$signed( -{ 2'b0,x458 }<<<3'd1 )+$signed( -{ 1'b0,x714 } )+$signed( { 1'b0,x203 }  )+$signed( { 1'b0,x459 }  )+$signed( { 1'b0,x715 }  )+$signed( -{ 2'b0,x474 }<<<3'd1 )+$signed( -{ 2'b0,x730 }<<<3'd1 )+$signed( { 2'b0,x475 } <<<3'd1 )+$signed( { 2'b0,x731 } <<<3'd1 )-$signed(11'd16);
assign y53=temp_y[53][11] ==1'b1 ? 5'd0 :  
        temp_y[53][8] ==1'b1 ? 5'd31 : 
        temp_y[53][2]==1'b1 ? temp_y[53][7:3]+1'b1 : temp_y[53][7:3];
assign temp_y[117] = 
+$signed( { 3'b0,x202 }<<<3'd2 )+$signed( -{ 2'b0,x458 }<<<3'd1 )+$signed( -{ 2'b0,x714 }<<<3'd1 )+$signed( { 2'b0,x203 } <<<3'd1 )+$signed( -{ 3'b0,x459 }<<<3'd2)+$signed( { 1'b0,x715 }  )+$signed( -{ 1'b0,x218 } )+$signed( { 1'b0,x730 }  )+$signed( -{ 2'b0,x219 }<<<3'd1 )+$signed( -{ 1'b0,x475 } )+$signed( { 2'b0,x731 } <<<3'd1 )+$signed(11'd24);
assign y117=temp_y[117][11] ==1'b1 ? 5'd0 :  
        temp_y[117][8] ==1'b1 ? 5'd31 : 
        temp_y[117][2]==1'b1 ? temp_y[117][7:3]+1'b1 : temp_y[117][7:3];
assign temp_y[181] = 
+$signed( { 2'b0,x202 } <<<3'd1 )+$signed( { 2'b0,x458 } <<<3'd1 )+$signed( { 1'b0,x714 }  )+$signed( { 2'b0,x203 } <<<3'd1 )+$signed( -{ 1'b0,x459 } )+$signed( { 1'b0,x715 }  )+$signed( -{ 2'b0,x218 }<<<3'd1 )+$signed( -{ 2'b0,x474 }<<<3'd1 )+$signed( -{ 1'b0,x730 } )+$signed( -{ 1'b0,x219 } )+$signed( -{ 1'b0,x475 } )+$signed( -{ 1'b0,x731 } )+$signed(11'd16);
assign y181=temp_y[181][11] ==1'b1 ? 5'd0 :  
        temp_y[181][8] ==1'b1 ? 5'd31 : 
        temp_y[181][2]==1'b1 ? temp_y[181][7:3]+1'b1 : temp_y[181][7:3];
assign temp_y[245] = 
+$signed( { 1'b0,x202 }  )+$signed( -{ 1'b0,x458 } )+$signed( { 1'b0,x203 }  )+$signed( -{ 1'b0,x459 } )+$signed( { 2'b0,x218 } <<<3'd1 )+$signed( -{ 1'b0,x474 } )+$signed( -{ 1'b0,x730 } )+$signed( { 2'b0,x219 } <<<3'd1 )+$signed( -{ 1'b0,x475 } )+$signed( -{ 2'b0,x731 }<<<3'd1 )+$signed(11'd40);
assign y245=temp_y[245][11] ==1'b1 ? 5'd0 :  
        temp_y[245][8] ==1'b1 ? 5'd31 : 
        temp_y[245][2]==1'b1 ? temp_y[245][7:3]+1'b1 : temp_y[245][7:3];
assign temp_y[309] = 
+$signed( -{ 1'b0,x202 } )+$signed( { 2'b0,x458 } <<<3'd1 )+$signed( -{ 1'b0,x714 } )+$signed( -{ 1'b0,x203 } )+$signed( { 2'b0,x459 } <<<3'd1 )+$signed( -{ 2'b0,x715 }<<<3'd1 )+$signed( -{ 1'b0,x218 } )+$signed( { 2'b0,x474 } <<<3'd1 )+$signed( -{ 1'b0,x730 } )+$signed( -{ 2'b0,x219 }<<<3'd1 )+$signed( { 3'b0,x475 }<<<3'd2 )+$signed( -{ 2'b0,x731 }<<<3'd1 )+$signed(11'd32);
assign y309=temp_y[309][11] ==1'b1 ? 5'd0 :  
        temp_y[309][8] ==1'b1 ? 5'd31 : 
        temp_y[309][2]==1'b1 ? temp_y[309][7:3]+1'b1 : temp_y[309][7:3];
assign temp_y[373] = 
+$signed( -{ 1'b0,x202 } )+$signed( -{ 2'b0,x458 }<<<3'd1 )+$signed( -{ 1'b0,x714 } )+$signed( { 1'b0,x203 }  )+$signed( { 2'b0,x459 } <<<3'd1 )+$signed( { 1'b0,x715 }  )+$signed( { 1'b0,x218 }  )+$signed( { 2'b0,x474 } <<<3'd1 )+$signed( { 2'b0,x730 } <<<3'd1 )+$signed( -{ 1'b0,x219 } )+$signed( -{ 2'b0,x475 }<<<3'd1 )+$signed( -{ 1'b0,x731 } )-$signed(11'd68);
assign y373=temp_y[373][11] ==1'b1 ? 5'd0 :  
        temp_y[373][8] ==1'b1 ? 5'd31 : 
        temp_y[373][2]==1'b1 ? temp_y[373][7:3]+1'b1 : temp_y[373][7:3];
assign temp_y[437] = 
+$signed( { 1'b0,x458 }  )+$signed( { 1'b0,x715 }  )+$signed( { 1'b0,x731 }  )-$signed(11'd108);
assign y437=temp_y[437][11] ==1'b1 ? 5'd0 :  
        temp_y[437][8] ==1'b1 ? 5'd31 : 
        temp_y[437][2]==1'b1 ? temp_y[437][7:3]+1'b1 : temp_y[437][7:3];
assign temp_y[501] = 
+$signed( -{ 2'b0,x202 }<<<3'd1 )+$signed( { 2'b0,x714 } <<<3'd1 )+$signed( -{ 2'b0,x203 }<<<3'd1 )+$signed( { 1'b0,x459 }  )+$signed( { 1'b0,x715 }  )+$signed( -{ 2'b0,x218 }<<<3'd1 )+$signed( { 1'b0,x474 }  )+$signed( { 1'b0,x730 }  )+$signed( -{ 1'b0,x219 } )+$signed(11'd64);
assign y501=temp_y[501][11] ==1'b1 ? 5'd0 :  
        temp_y[501][8] ==1'b1 ? 5'd31 : 
        temp_y[501][2]==1'b1 ? temp_y[501][7:3]+1'b1 : temp_y[501][7:3];
assign temp_y[565] = 
+$signed( -{ 2'b0,x202 }<<<3'd1 )+$signed( -{ 1'b0,x458 } )+$signed( -{ 3'b0,x203 }<<<3'd2)+$signed( { 1'b0,x218 }  )+$signed( { 1'b0,x474 }  )+$signed( { 3'b0,x219 }<<<3'd2 )+$signed(11'd16);
assign y565=temp_y[565][11] ==1'b1 ? 5'd0 :  
        temp_y[565][8] ==1'b1 ? 5'd31 : 
        temp_y[565][2]==1'b1 ? temp_y[565][7:3]+1'b1 : temp_y[565][7:3];
assign temp_y[629] = 
+$signed( { 2'b0,x458 } <<<3'd1 )+$signed( { 2'b0,x714 } <<<3'd1 )+$signed( -{ 1'b0,x203 } )+$signed( -{ 2'b0,x459 }<<<3'd1 )+$signed( -{ 2'b0,x715 }<<<3'd1 )+$signed( { 2'b0,x474 } <<<3'd1 )+$signed( { 1'b0,x730 }  )+$signed( -{ 2'b0,x475 }<<<3'd1 )-$signed(11'd8);
assign y629=temp_y[629][11] ==1'b1 ? 5'd0 :  
        temp_y[629][8] ==1'b1 ? 5'd31 : 
        temp_y[629][2]==1'b1 ? temp_y[629][7:3]+1'b1 : temp_y[629][7:3];
assign temp_y[54] = 
+$signed( -{ 2'b0,x460 }<<<3'd1 )+$signed( -{ 1'b0,x716 } )+$signed( { 1'b0,x205 }  )+$signed( { 1'b0,x461 }  )+$signed( { 1'b0,x717 }  )+$signed( -{ 2'b0,x476 }<<<3'd1 )+$signed( -{ 2'b0,x732 }<<<3'd1 )+$signed( { 2'b0,x477 } <<<3'd1 )+$signed( { 2'b0,x733 } <<<3'd1 )-$signed(11'd16);
assign y54=temp_y[54][11] ==1'b1 ? 5'd0 :  
        temp_y[54][8] ==1'b1 ? 5'd31 : 
        temp_y[54][2]==1'b1 ? temp_y[54][7:3]+1'b1 : temp_y[54][7:3];
assign temp_y[118] = 
+$signed( { 3'b0,x204 }<<<3'd2 )+$signed( -{ 2'b0,x460 }<<<3'd1 )+$signed( -{ 2'b0,x716 }<<<3'd1 )+$signed( { 2'b0,x205 } <<<3'd1 )+$signed( -{ 3'b0,x461 }<<<3'd2)+$signed( { 1'b0,x717 }  )+$signed( -{ 1'b0,x220 } )+$signed( { 1'b0,x732 }  )+$signed( -{ 2'b0,x221 }<<<3'd1 )+$signed( -{ 1'b0,x477 } )+$signed( { 2'b0,x733 } <<<3'd1 )+$signed(11'd24);
assign y118=temp_y[118][11] ==1'b1 ? 5'd0 :  
        temp_y[118][8] ==1'b1 ? 5'd31 : 
        temp_y[118][2]==1'b1 ? temp_y[118][7:3]+1'b1 : temp_y[118][7:3];
assign temp_y[182] = 
+$signed( { 2'b0,x204 } <<<3'd1 )+$signed( { 2'b0,x460 } <<<3'd1 )+$signed( { 1'b0,x716 }  )+$signed( { 2'b0,x205 } <<<3'd1 )+$signed( -{ 1'b0,x461 } )+$signed( { 1'b0,x717 }  )+$signed( -{ 2'b0,x220 }<<<3'd1 )+$signed( -{ 2'b0,x476 }<<<3'd1 )+$signed( -{ 1'b0,x732 } )+$signed( -{ 1'b0,x221 } )+$signed( -{ 1'b0,x477 } )+$signed( -{ 1'b0,x733 } )+$signed(11'd16);
assign y182=temp_y[182][11] ==1'b1 ? 5'd0 :  
        temp_y[182][8] ==1'b1 ? 5'd31 : 
        temp_y[182][2]==1'b1 ? temp_y[182][7:3]+1'b1 : temp_y[182][7:3];
assign temp_y[246] = 
+$signed( { 1'b0,x204 }  )+$signed( -{ 1'b0,x460 } )+$signed( { 1'b0,x205 }  )+$signed( -{ 1'b0,x461 } )+$signed( { 2'b0,x220 } <<<3'd1 )+$signed( -{ 1'b0,x476 } )+$signed( -{ 1'b0,x732 } )+$signed( { 2'b0,x221 } <<<3'd1 )+$signed( -{ 1'b0,x477 } )+$signed( -{ 2'b0,x733 }<<<3'd1 )+$signed(11'd40);
assign y246=temp_y[246][11] ==1'b1 ? 5'd0 :  
        temp_y[246][8] ==1'b1 ? 5'd31 : 
        temp_y[246][2]==1'b1 ? temp_y[246][7:3]+1'b1 : temp_y[246][7:3];
assign temp_y[310] = 
+$signed( -{ 1'b0,x204 } )+$signed( { 2'b0,x460 } <<<3'd1 )+$signed( -{ 1'b0,x716 } )+$signed( -{ 1'b0,x205 } )+$signed( { 2'b0,x461 } <<<3'd1 )+$signed( -{ 2'b0,x717 }<<<3'd1 )+$signed( -{ 1'b0,x220 } )+$signed( { 2'b0,x476 } <<<3'd1 )+$signed( -{ 1'b0,x732 } )+$signed( -{ 2'b0,x221 }<<<3'd1 )+$signed( { 3'b0,x477 }<<<3'd2 )+$signed( -{ 2'b0,x733 }<<<3'd1 )+$signed(11'd32);
assign y310=temp_y[310][11] ==1'b1 ? 5'd0 :  
        temp_y[310][8] ==1'b1 ? 5'd31 : 
        temp_y[310][2]==1'b1 ? temp_y[310][7:3]+1'b1 : temp_y[310][7:3];
assign temp_y[374] = 
+$signed( -{ 1'b0,x204 } )+$signed( -{ 2'b0,x460 }<<<3'd1 )+$signed( -{ 1'b0,x716 } )+$signed( { 1'b0,x205 }  )+$signed( { 2'b0,x461 } <<<3'd1 )+$signed( { 1'b0,x717 }  )+$signed( { 1'b0,x220 }  )+$signed( { 2'b0,x476 } <<<3'd1 )+$signed( { 2'b0,x732 } <<<3'd1 )+$signed( -{ 1'b0,x221 } )+$signed( -{ 2'b0,x477 }<<<3'd1 )+$signed( -{ 1'b0,x733 } )-$signed(11'd68);
assign y374=temp_y[374][11] ==1'b1 ? 5'd0 :  
        temp_y[374][8] ==1'b1 ? 5'd31 : 
        temp_y[374][2]==1'b1 ? temp_y[374][7:3]+1'b1 : temp_y[374][7:3];
assign temp_y[438] = 
+$signed( { 1'b0,x460 }  )+$signed( { 1'b0,x717 }  )+$signed( { 1'b0,x733 }  )-$signed(11'd108);
assign y438=temp_y[438][11] ==1'b1 ? 5'd0 :  
        temp_y[438][8] ==1'b1 ? 5'd31 : 
        temp_y[438][2]==1'b1 ? temp_y[438][7:3]+1'b1 : temp_y[438][7:3];
assign temp_y[502] = 
+$signed( -{ 2'b0,x204 }<<<3'd1 )+$signed( { 2'b0,x716 } <<<3'd1 )+$signed( -{ 2'b0,x205 }<<<3'd1 )+$signed( { 1'b0,x461 }  )+$signed( { 1'b0,x717 }  )+$signed( -{ 2'b0,x220 }<<<3'd1 )+$signed( { 1'b0,x476 }  )+$signed( { 1'b0,x732 }  )+$signed( -{ 1'b0,x221 } )+$signed(11'd64);
assign y502=temp_y[502][11] ==1'b1 ? 5'd0 :  
        temp_y[502][8] ==1'b1 ? 5'd31 : 
        temp_y[502][2]==1'b1 ? temp_y[502][7:3]+1'b1 : temp_y[502][7:3];
assign temp_y[566] = 
+$signed( -{ 2'b0,x204 }<<<3'd1 )+$signed( -{ 1'b0,x460 } )+$signed( -{ 3'b0,x205 }<<<3'd2)+$signed( { 1'b0,x220 }  )+$signed( { 1'b0,x476 }  )+$signed( { 3'b0,x221 }<<<3'd2 )+$signed(11'd16);
assign y566=temp_y[566][11] ==1'b1 ? 5'd0 :  
        temp_y[566][8] ==1'b1 ? 5'd31 : 
        temp_y[566][2]==1'b1 ? temp_y[566][7:3]+1'b1 : temp_y[566][7:3];
assign temp_y[630] = 
+$signed( { 2'b0,x460 } <<<3'd1 )+$signed( { 2'b0,x716 } <<<3'd1 )+$signed( -{ 1'b0,x205 } )+$signed( -{ 2'b0,x461 }<<<3'd1 )+$signed( -{ 2'b0,x717 }<<<3'd1 )+$signed( { 2'b0,x476 } <<<3'd1 )+$signed( { 1'b0,x732 }  )+$signed( -{ 2'b0,x477 }<<<3'd1 )-$signed(11'd8);
assign y630=temp_y[630][11] ==1'b1 ? 5'd0 :  
        temp_y[630][8] ==1'b1 ? 5'd31 : 
        temp_y[630][2]==1'b1 ? temp_y[630][7:3]+1'b1 : temp_y[630][7:3];
assign temp_y[55] = 
+$signed( -{ 2'b0,x462 }<<<3'd1 )+$signed( -{ 1'b0,x718 } )+$signed( { 1'b0,x207 }  )+$signed( { 1'b0,x463 }  )+$signed( { 1'b0,x719 }  )+$signed( -{ 2'b0,x478 }<<<3'd1 )+$signed( -{ 2'b0,x734 }<<<3'd1 )+$signed( { 2'b0,x479 } <<<3'd1 )+$signed( { 2'b0,x735 } <<<3'd1 )-$signed(11'd16);
assign y55=temp_y[55][11] ==1'b1 ? 5'd0 :  
        temp_y[55][8] ==1'b1 ? 5'd31 : 
        temp_y[55][2]==1'b1 ? temp_y[55][7:3]+1'b1 : temp_y[55][7:3];
assign temp_y[119] = 
+$signed( { 3'b0,x206 }<<<3'd2 )+$signed( -{ 2'b0,x462 }<<<3'd1 )+$signed( -{ 2'b0,x718 }<<<3'd1 )+$signed( { 2'b0,x207 } <<<3'd1 )+$signed( -{ 3'b0,x463 }<<<3'd2)+$signed( { 1'b0,x719 }  )+$signed( -{ 1'b0,x222 } )+$signed( { 1'b0,x734 }  )+$signed( -{ 2'b0,x223 }<<<3'd1 )+$signed( -{ 1'b0,x479 } )+$signed( { 2'b0,x735 } <<<3'd1 )+$signed(11'd24);
assign y119=temp_y[119][11] ==1'b1 ? 5'd0 :  
        temp_y[119][8] ==1'b1 ? 5'd31 : 
        temp_y[119][2]==1'b1 ? temp_y[119][7:3]+1'b1 : temp_y[119][7:3];
assign temp_y[183] = 
+$signed( { 2'b0,x206 } <<<3'd1 )+$signed( { 2'b0,x462 } <<<3'd1 )+$signed( { 1'b0,x718 }  )+$signed( { 2'b0,x207 } <<<3'd1 )+$signed( -{ 1'b0,x463 } )+$signed( { 1'b0,x719 }  )+$signed( -{ 2'b0,x222 }<<<3'd1 )+$signed( -{ 2'b0,x478 }<<<3'd1 )+$signed( -{ 1'b0,x734 } )+$signed( -{ 1'b0,x223 } )+$signed( -{ 1'b0,x479 } )+$signed( -{ 1'b0,x735 } )+$signed(11'd16);
assign y183=temp_y[183][11] ==1'b1 ? 5'd0 :  
        temp_y[183][8] ==1'b1 ? 5'd31 : 
        temp_y[183][2]==1'b1 ? temp_y[183][7:3]+1'b1 : temp_y[183][7:3];
assign temp_y[247] = 
+$signed( { 1'b0,x206 }  )+$signed( -{ 1'b0,x462 } )+$signed( { 1'b0,x207 }  )+$signed( -{ 1'b0,x463 } )+$signed( { 2'b0,x222 } <<<3'd1 )+$signed( -{ 1'b0,x478 } )+$signed( -{ 1'b0,x734 } )+$signed( { 2'b0,x223 } <<<3'd1 )+$signed( -{ 1'b0,x479 } )+$signed( -{ 2'b0,x735 }<<<3'd1 )+$signed(11'd40);
assign y247=temp_y[247][11] ==1'b1 ? 5'd0 :  
        temp_y[247][8] ==1'b1 ? 5'd31 : 
        temp_y[247][2]==1'b1 ? temp_y[247][7:3]+1'b1 : temp_y[247][7:3];
assign temp_y[311] = 
+$signed( -{ 1'b0,x206 } )+$signed( { 2'b0,x462 } <<<3'd1 )+$signed( -{ 1'b0,x718 } )+$signed( -{ 1'b0,x207 } )+$signed( { 2'b0,x463 } <<<3'd1 )+$signed( -{ 2'b0,x719 }<<<3'd1 )+$signed( -{ 1'b0,x222 } )+$signed( { 2'b0,x478 } <<<3'd1 )+$signed( -{ 1'b0,x734 } )+$signed( -{ 2'b0,x223 }<<<3'd1 )+$signed( { 3'b0,x479 }<<<3'd2 )+$signed( -{ 2'b0,x735 }<<<3'd1 )+$signed(11'd32);
assign y311=temp_y[311][11] ==1'b1 ? 5'd0 :  
        temp_y[311][8] ==1'b1 ? 5'd31 : 
        temp_y[311][2]==1'b1 ? temp_y[311][7:3]+1'b1 : temp_y[311][7:3];
assign temp_y[375] = 
+$signed( -{ 1'b0,x206 } )+$signed( -{ 2'b0,x462 }<<<3'd1 )+$signed( -{ 1'b0,x718 } )+$signed( { 1'b0,x207 }  )+$signed( { 2'b0,x463 } <<<3'd1 )+$signed( { 1'b0,x719 }  )+$signed( { 1'b0,x222 }  )+$signed( { 2'b0,x478 } <<<3'd1 )+$signed( { 2'b0,x734 } <<<3'd1 )+$signed( -{ 1'b0,x223 } )+$signed( -{ 2'b0,x479 }<<<3'd1 )+$signed( -{ 1'b0,x735 } )-$signed(11'd68);
assign y375=temp_y[375][11] ==1'b1 ? 5'd0 :  
        temp_y[375][8] ==1'b1 ? 5'd31 : 
        temp_y[375][2]==1'b1 ? temp_y[375][7:3]+1'b1 : temp_y[375][7:3];
assign temp_y[439] = 
+$signed( { 1'b0,x462 }  )+$signed( { 1'b0,x719 }  )+$signed( { 1'b0,x735 }  )-$signed(11'd108);
assign y439=temp_y[439][11] ==1'b1 ? 5'd0 :  
        temp_y[439][8] ==1'b1 ? 5'd31 : 
        temp_y[439][2]==1'b1 ? temp_y[439][7:3]+1'b1 : temp_y[439][7:3];
assign temp_y[503] = 
+$signed( -{ 2'b0,x206 }<<<3'd1 )+$signed( { 2'b0,x718 } <<<3'd1 )+$signed( -{ 2'b0,x207 }<<<3'd1 )+$signed( { 1'b0,x463 }  )+$signed( { 1'b0,x719 }  )+$signed( -{ 2'b0,x222 }<<<3'd1 )+$signed( { 1'b0,x478 }  )+$signed( { 1'b0,x734 }  )+$signed( -{ 1'b0,x223 } )+$signed(11'd64);
assign y503=temp_y[503][11] ==1'b1 ? 5'd0 :  
        temp_y[503][8] ==1'b1 ? 5'd31 : 
        temp_y[503][2]==1'b1 ? temp_y[503][7:3]+1'b1 : temp_y[503][7:3];
assign temp_y[567] = 
+$signed( -{ 2'b0,x206 }<<<3'd1 )+$signed( -{ 1'b0,x462 } )+$signed( -{ 3'b0,x207 }<<<3'd2)+$signed( { 1'b0,x222 }  )+$signed( { 1'b0,x478 }  )+$signed( { 3'b0,x223 }<<<3'd2 )+$signed(11'd16);
assign y567=temp_y[567][11] ==1'b1 ? 5'd0 :  
        temp_y[567][8] ==1'b1 ? 5'd31 : 
        temp_y[567][2]==1'b1 ? temp_y[567][7:3]+1'b1 : temp_y[567][7:3];
assign temp_y[631] = 
+$signed( { 2'b0,x462 } <<<3'd1 )+$signed( { 2'b0,x718 } <<<3'd1 )+$signed( -{ 1'b0,x207 } )+$signed( -{ 2'b0,x463 }<<<3'd1 )+$signed( -{ 2'b0,x719 }<<<3'd1 )+$signed( { 2'b0,x478 } <<<3'd1 )+$signed( { 1'b0,x734 }  )+$signed( -{ 2'b0,x479 }<<<3'd1 )-$signed(11'd8);
assign y631=temp_y[631][11] ==1'b1 ? 5'd0 :  
        temp_y[631][8] ==1'b1 ? 5'd31 : 
        temp_y[631][2]==1'b1 ? temp_y[631][7:3]+1'b1 : temp_y[631][7:3];
assign temp_y[56] = 
+$signed( -{ 2'b0,x480 }<<<3'd1 )+$signed( -{ 1'b0,x736 } )+$signed( { 1'b0,x225 }  )+$signed( { 1'b0,x481 }  )+$signed( { 1'b0,x737 }  )+$signed( -{ 2'b0,x496 }<<<3'd1 )+$signed( -{ 2'b0,x752 }<<<3'd1 )+$signed( { 2'b0,x497 } <<<3'd1 )+$signed( { 2'b0,x753 } <<<3'd1 )-$signed(11'd16);
assign y56=temp_y[56][11] ==1'b1 ? 5'd0 :  
        temp_y[56][8] ==1'b1 ? 5'd31 : 
        temp_y[56][2]==1'b1 ? temp_y[56][7:3]+1'b1 : temp_y[56][7:3];
assign temp_y[120] = 
+$signed( { 3'b0,x224 }<<<3'd2 )+$signed( -{ 2'b0,x480 }<<<3'd1 )+$signed( -{ 2'b0,x736 }<<<3'd1 )+$signed( { 2'b0,x225 } <<<3'd1 )+$signed( -{ 3'b0,x481 }<<<3'd2)+$signed( { 1'b0,x737 }  )+$signed( -{ 1'b0,x240 } )+$signed( { 1'b0,x752 }  )+$signed( -{ 2'b0,x241 }<<<3'd1 )+$signed( -{ 1'b0,x497 } )+$signed( { 2'b0,x753 } <<<3'd1 )+$signed(11'd24);
assign y120=temp_y[120][11] ==1'b1 ? 5'd0 :  
        temp_y[120][8] ==1'b1 ? 5'd31 : 
        temp_y[120][2]==1'b1 ? temp_y[120][7:3]+1'b1 : temp_y[120][7:3];
assign temp_y[184] = 
+$signed( { 2'b0,x224 } <<<3'd1 )+$signed( { 2'b0,x480 } <<<3'd1 )+$signed( { 1'b0,x736 }  )+$signed( { 2'b0,x225 } <<<3'd1 )+$signed( -{ 1'b0,x481 } )+$signed( { 1'b0,x737 }  )+$signed( -{ 2'b0,x240 }<<<3'd1 )+$signed( -{ 2'b0,x496 }<<<3'd1 )+$signed( -{ 1'b0,x752 } )+$signed( -{ 1'b0,x241 } )+$signed( -{ 1'b0,x497 } )+$signed( -{ 1'b0,x753 } )+$signed(11'd16);
assign y184=temp_y[184][11] ==1'b1 ? 5'd0 :  
        temp_y[184][8] ==1'b1 ? 5'd31 : 
        temp_y[184][2]==1'b1 ? temp_y[184][7:3]+1'b1 : temp_y[184][7:3];
assign temp_y[248] = 
+$signed( { 1'b0,x224 }  )+$signed( -{ 1'b0,x480 } )+$signed( { 1'b0,x225 }  )+$signed( -{ 1'b0,x481 } )+$signed( { 2'b0,x240 } <<<3'd1 )+$signed( -{ 1'b0,x496 } )+$signed( -{ 1'b0,x752 } )+$signed( { 2'b0,x241 } <<<3'd1 )+$signed( -{ 1'b0,x497 } )+$signed( -{ 2'b0,x753 }<<<3'd1 )+$signed(11'd40);
assign y248=temp_y[248][11] ==1'b1 ? 5'd0 :  
        temp_y[248][8] ==1'b1 ? 5'd31 : 
        temp_y[248][2]==1'b1 ? temp_y[248][7:3]+1'b1 : temp_y[248][7:3];
assign temp_y[312] = 
+$signed( -{ 1'b0,x224 } )+$signed( { 2'b0,x480 } <<<3'd1 )+$signed( -{ 1'b0,x736 } )+$signed( -{ 1'b0,x225 } )+$signed( { 2'b0,x481 } <<<3'd1 )+$signed( -{ 2'b0,x737 }<<<3'd1 )+$signed( -{ 1'b0,x240 } )+$signed( { 2'b0,x496 } <<<3'd1 )+$signed( -{ 1'b0,x752 } )+$signed( -{ 2'b0,x241 }<<<3'd1 )+$signed( { 3'b0,x497 }<<<3'd2 )+$signed( -{ 2'b0,x753 }<<<3'd1 )+$signed(11'd32);
assign y312=temp_y[312][11] ==1'b1 ? 5'd0 :  
        temp_y[312][8] ==1'b1 ? 5'd31 : 
        temp_y[312][2]==1'b1 ? temp_y[312][7:3]+1'b1 : temp_y[312][7:3];
assign temp_y[376] = 
+$signed( -{ 1'b0,x224 } )+$signed( -{ 2'b0,x480 }<<<3'd1 )+$signed( -{ 1'b0,x736 } )+$signed( { 1'b0,x225 }  )+$signed( { 2'b0,x481 } <<<3'd1 )+$signed( { 1'b0,x737 }  )+$signed( { 1'b0,x240 }  )+$signed( { 2'b0,x496 } <<<3'd1 )+$signed( { 2'b0,x752 } <<<3'd1 )+$signed( -{ 1'b0,x241 } )+$signed( -{ 2'b0,x497 }<<<3'd1 )+$signed( -{ 1'b0,x753 } )-$signed(11'd68);
assign y376=temp_y[376][11] ==1'b1 ? 5'd0 :  
        temp_y[376][8] ==1'b1 ? 5'd31 : 
        temp_y[376][2]==1'b1 ? temp_y[376][7:3]+1'b1 : temp_y[376][7:3];
assign temp_y[440] = 
+$signed( { 1'b0,x480 }  )+$signed( { 1'b0,x737 }  )+$signed( { 1'b0,x753 }  )-$signed(11'd108);
assign y440=temp_y[440][11] ==1'b1 ? 5'd0 :  
        temp_y[440][8] ==1'b1 ? 5'd31 : 
        temp_y[440][2]==1'b1 ? temp_y[440][7:3]+1'b1 : temp_y[440][7:3];
assign temp_y[504] = 
+$signed( -{ 2'b0,x224 }<<<3'd1 )+$signed( { 2'b0,x736 } <<<3'd1 )+$signed( -{ 2'b0,x225 }<<<3'd1 )+$signed( { 1'b0,x481 }  )+$signed( { 1'b0,x737 }  )+$signed( -{ 2'b0,x240 }<<<3'd1 )+$signed( { 1'b0,x496 }  )+$signed( { 1'b0,x752 }  )+$signed( -{ 1'b0,x241 } )+$signed(11'd64);
assign y504=temp_y[504][11] ==1'b1 ? 5'd0 :  
        temp_y[504][8] ==1'b1 ? 5'd31 : 
        temp_y[504][2]==1'b1 ? temp_y[504][7:3]+1'b1 : temp_y[504][7:3];
assign temp_y[568] = 
+$signed( -{ 2'b0,x224 }<<<3'd1 )+$signed( -{ 1'b0,x480 } )+$signed( -{ 3'b0,x225 }<<<3'd2)+$signed( { 1'b0,x240 }  )+$signed( { 1'b0,x496 }  )+$signed( { 3'b0,x241 }<<<3'd2 )+$signed(11'd16);
assign y568=temp_y[568][11] ==1'b1 ? 5'd0 :  
        temp_y[568][8] ==1'b1 ? 5'd31 : 
        temp_y[568][2]==1'b1 ? temp_y[568][7:3]+1'b1 : temp_y[568][7:3];
assign temp_y[632] = 
+$signed( { 2'b0,x480 } <<<3'd1 )+$signed( { 2'b0,x736 } <<<3'd1 )+$signed( -{ 1'b0,x225 } )+$signed( -{ 2'b0,x481 }<<<3'd1 )+$signed( -{ 2'b0,x737 }<<<3'd1 )+$signed( { 2'b0,x496 } <<<3'd1 )+$signed( { 1'b0,x752 }  )+$signed( -{ 2'b0,x497 }<<<3'd1 )-$signed(11'd8);
assign y632=temp_y[632][11] ==1'b1 ? 5'd0 :  
        temp_y[632][8] ==1'b1 ? 5'd31 : 
        temp_y[632][2]==1'b1 ? temp_y[632][7:3]+1'b1 : temp_y[632][7:3];
assign temp_y[57] = 
+$signed( -{ 2'b0,x482 }<<<3'd1 )+$signed( -{ 1'b0,x738 } )+$signed( { 1'b0,x227 }  )+$signed( { 1'b0,x483 }  )+$signed( { 1'b0,x739 }  )+$signed( -{ 2'b0,x498 }<<<3'd1 )+$signed( -{ 2'b0,x754 }<<<3'd1 )+$signed( { 2'b0,x499 } <<<3'd1 )+$signed( { 2'b0,x755 } <<<3'd1 )-$signed(11'd16);
assign y57=temp_y[57][11] ==1'b1 ? 5'd0 :  
        temp_y[57][8] ==1'b1 ? 5'd31 : 
        temp_y[57][2]==1'b1 ? temp_y[57][7:3]+1'b1 : temp_y[57][7:3];
assign temp_y[121] = 
+$signed( { 3'b0,x226 }<<<3'd2 )+$signed( -{ 2'b0,x482 }<<<3'd1 )+$signed( -{ 2'b0,x738 }<<<3'd1 )+$signed( { 2'b0,x227 } <<<3'd1 )+$signed( -{ 3'b0,x483 }<<<3'd2)+$signed( { 1'b0,x739 }  )+$signed( -{ 1'b0,x242 } )+$signed( { 1'b0,x754 }  )+$signed( -{ 2'b0,x243 }<<<3'd1 )+$signed( -{ 1'b0,x499 } )+$signed( { 2'b0,x755 } <<<3'd1 )+$signed(11'd24);
assign y121=temp_y[121][11] ==1'b1 ? 5'd0 :  
        temp_y[121][8] ==1'b1 ? 5'd31 : 
        temp_y[121][2]==1'b1 ? temp_y[121][7:3]+1'b1 : temp_y[121][7:3];
assign temp_y[185] = 
+$signed( { 2'b0,x226 } <<<3'd1 )+$signed( { 2'b0,x482 } <<<3'd1 )+$signed( { 1'b0,x738 }  )+$signed( { 2'b0,x227 } <<<3'd1 )+$signed( -{ 1'b0,x483 } )+$signed( { 1'b0,x739 }  )+$signed( -{ 2'b0,x242 }<<<3'd1 )+$signed( -{ 2'b0,x498 }<<<3'd1 )+$signed( -{ 1'b0,x754 } )+$signed( -{ 1'b0,x243 } )+$signed( -{ 1'b0,x499 } )+$signed( -{ 1'b0,x755 } )+$signed(11'd16);
assign y185=temp_y[185][11] ==1'b1 ? 5'd0 :  
        temp_y[185][8] ==1'b1 ? 5'd31 : 
        temp_y[185][2]==1'b1 ? temp_y[185][7:3]+1'b1 : temp_y[185][7:3];
assign temp_y[249] = 
+$signed( { 1'b0,x226 }  )+$signed( -{ 1'b0,x482 } )+$signed( { 1'b0,x227 }  )+$signed( -{ 1'b0,x483 } )+$signed( { 2'b0,x242 } <<<3'd1 )+$signed( -{ 1'b0,x498 } )+$signed( -{ 1'b0,x754 } )+$signed( { 2'b0,x243 } <<<3'd1 )+$signed( -{ 1'b0,x499 } )+$signed( -{ 2'b0,x755 }<<<3'd1 )+$signed(11'd40);
assign y249=temp_y[249][11] ==1'b1 ? 5'd0 :  
        temp_y[249][8] ==1'b1 ? 5'd31 : 
        temp_y[249][2]==1'b1 ? temp_y[249][7:3]+1'b1 : temp_y[249][7:3];
assign temp_y[313] = 
+$signed( -{ 1'b0,x226 } )+$signed( { 2'b0,x482 } <<<3'd1 )+$signed( -{ 1'b0,x738 } )+$signed( -{ 1'b0,x227 } )+$signed( { 2'b0,x483 } <<<3'd1 )+$signed( -{ 2'b0,x739 }<<<3'd1 )+$signed( -{ 1'b0,x242 } )+$signed( { 2'b0,x498 } <<<3'd1 )+$signed( -{ 1'b0,x754 } )+$signed( -{ 2'b0,x243 }<<<3'd1 )+$signed( { 3'b0,x499 }<<<3'd2 )+$signed( -{ 2'b0,x755 }<<<3'd1 )+$signed(11'd32);
assign y313=temp_y[313][11] ==1'b1 ? 5'd0 :  
        temp_y[313][8] ==1'b1 ? 5'd31 : 
        temp_y[313][2]==1'b1 ? temp_y[313][7:3]+1'b1 : temp_y[313][7:3];
assign temp_y[377] = 
+$signed( -{ 1'b0,x226 } )+$signed( -{ 2'b0,x482 }<<<3'd1 )+$signed( -{ 1'b0,x738 } )+$signed( { 1'b0,x227 }  )+$signed( { 2'b0,x483 } <<<3'd1 )+$signed( { 1'b0,x739 }  )+$signed( { 1'b0,x242 }  )+$signed( { 2'b0,x498 } <<<3'd1 )+$signed( { 2'b0,x754 } <<<3'd1 )+$signed( -{ 1'b0,x243 } )+$signed( -{ 2'b0,x499 }<<<3'd1 )+$signed( -{ 1'b0,x755 } )-$signed(11'd68);
assign y377=temp_y[377][11] ==1'b1 ? 5'd0 :  
        temp_y[377][8] ==1'b1 ? 5'd31 : 
        temp_y[377][2]==1'b1 ? temp_y[377][7:3]+1'b1 : temp_y[377][7:3];
assign temp_y[441] = 
+$signed( { 1'b0,x482 }  )+$signed( { 1'b0,x739 }  )+$signed( { 1'b0,x755 }  )-$signed(11'd108);
assign y441=temp_y[441][11] ==1'b1 ? 5'd0 :  
        temp_y[441][8] ==1'b1 ? 5'd31 : 
        temp_y[441][2]==1'b1 ? temp_y[441][7:3]+1'b1 : temp_y[441][7:3];
assign temp_y[505] = 
+$signed( -{ 2'b0,x226 }<<<3'd1 )+$signed( { 2'b0,x738 } <<<3'd1 )+$signed( -{ 2'b0,x227 }<<<3'd1 )+$signed( { 1'b0,x483 }  )+$signed( { 1'b0,x739 }  )+$signed( -{ 2'b0,x242 }<<<3'd1 )+$signed( { 1'b0,x498 }  )+$signed( { 1'b0,x754 }  )+$signed( -{ 1'b0,x243 } )+$signed(11'd64);
assign y505=temp_y[505][11] ==1'b1 ? 5'd0 :  
        temp_y[505][8] ==1'b1 ? 5'd31 : 
        temp_y[505][2]==1'b1 ? temp_y[505][7:3]+1'b1 : temp_y[505][7:3];
assign temp_y[569] = 
+$signed( -{ 2'b0,x226 }<<<3'd1 )+$signed( -{ 1'b0,x482 } )+$signed( -{ 3'b0,x227 }<<<3'd2)+$signed( { 1'b0,x242 }  )+$signed( { 1'b0,x498 }  )+$signed( { 3'b0,x243 }<<<3'd2 )+$signed(11'd16);
assign y569=temp_y[569][11] ==1'b1 ? 5'd0 :  
        temp_y[569][8] ==1'b1 ? 5'd31 : 
        temp_y[569][2]==1'b1 ? temp_y[569][7:3]+1'b1 : temp_y[569][7:3];
assign temp_y[633] = 
+$signed( { 2'b0,x482 } <<<3'd1 )+$signed( { 2'b0,x738 } <<<3'd1 )+$signed( -{ 1'b0,x227 } )+$signed( -{ 2'b0,x483 }<<<3'd1 )+$signed( -{ 2'b0,x739 }<<<3'd1 )+$signed( { 2'b0,x498 } <<<3'd1 )+$signed( { 1'b0,x754 }  )+$signed( -{ 2'b0,x499 }<<<3'd1 )-$signed(11'd8);
assign y633=temp_y[633][11] ==1'b1 ? 5'd0 :  
        temp_y[633][8] ==1'b1 ? 5'd31 : 
        temp_y[633][2]==1'b1 ? temp_y[633][7:3]+1'b1 : temp_y[633][7:3];
assign temp_y[58] = 
+$signed( -{ 2'b0,x484 }<<<3'd1 )+$signed( -{ 1'b0,x740 } )+$signed( { 1'b0,x229 }  )+$signed( { 1'b0,x485 }  )+$signed( { 1'b0,x741 }  )+$signed( -{ 2'b0,x500 }<<<3'd1 )+$signed( -{ 2'b0,x756 }<<<3'd1 )+$signed( { 2'b0,x501 } <<<3'd1 )+$signed( { 2'b0,x757 } <<<3'd1 )-$signed(11'd16);
assign y58=temp_y[58][11] ==1'b1 ? 5'd0 :  
        temp_y[58][8] ==1'b1 ? 5'd31 : 
        temp_y[58][2]==1'b1 ? temp_y[58][7:3]+1'b1 : temp_y[58][7:3];
assign temp_y[122] = 
+$signed( { 3'b0,x228 }<<<3'd2 )+$signed( -{ 2'b0,x484 }<<<3'd1 )+$signed( -{ 2'b0,x740 }<<<3'd1 )+$signed( { 2'b0,x229 } <<<3'd1 )+$signed( -{ 3'b0,x485 }<<<3'd2)+$signed( { 1'b0,x741 }  )+$signed( -{ 1'b0,x244 } )+$signed( { 1'b0,x756 }  )+$signed( -{ 2'b0,x245 }<<<3'd1 )+$signed( -{ 1'b0,x501 } )+$signed( { 2'b0,x757 } <<<3'd1 )+$signed(11'd24);
assign y122=temp_y[122][11] ==1'b1 ? 5'd0 :  
        temp_y[122][8] ==1'b1 ? 5'd31 : 
        temp_y[122][2]==1'b1 ? temp_y[122][7:3]+1'b1 : temp_y[122][7:3];
assign temp_y[186] = 
+$signed( { 2'b0,x228 } <<<3'd1 )+$signed( { 2'b0,x484 } <<<3'd1 )+$signed( { 1'b0,x740 }  )+$signed( { 2'b0,x229 } <<<3'd1 )+$signed( -{ 1'b0,x485 } )+$signed( { 1'b0,x741 }  )+$signed( -{ 2'b0,x244 }<<<3'd1 )+$signed( -{ 2'b0,x500 }<<<3'd1 )+$signed( -{ 1'b0,x756 } )+$signed( -{ 1'b0,x245 } )+$signed( -{ 1'b0,x501 } )+$signed( -{ 1'b0,x757 } )+$signed(11'd16);
assign y186=temp_y[186][11] ==1'b1 ? 5'd0 :  
        temp_y[186][8] ==1'b1 ? 5'd31 : 
        temp_y[186][2]==1'b1 ? temp_y[186][7:3]+1'b1 : temp_y[186][7:3];
assign temp_y[250] = 
+$signed( { 1'b0,x228 }  )+$signed( -{ 1'b0,x484 } )+$signed( { 1'b0,x229 }  )+$signed( -{ 1'b0,x485 } )+$signed( { 2'b0,x244 } <<<3'd1 )+$signed( -{ 1'b0,x500 } )+$signed( -{ 1'b0,x756 } )+$signed( { 2'b0,x245 } <<<3'd1 )+$signed( -{ 1'b0,x501 } )+$signed( -{ 2'b0,x757 }<<<3'd1 )+$signed(11'd40);
assign y250=temp_y[250][11] ==1'b1 ? 5'd0 :  
        temp_y[250][8] ==1'b1 ? 5'd31 : 
        temp_y[250][2]==1'b1 ? temp_y[250][7:3]+1'b1 : temp_y[250][7:3];
assign temp_y[314] = 
+$signed( -{ 1'b0,x228 } )+$signed( { 2'b0,x484 } <<<3'd1 )+$signed( -{ 1'b0,x740 } )+$signed( -{ 1'b0,x229 } )+$signed( { 2'b0,x485 } <<<3'd1 )+$signed( -{ 2'b0,x741 }<<<3'd1 )+$signed( -{ 1'b0,x244 } )+$signed( { 2'b0,x500 } <<<3'd1 )+$signed( -{ 1'b0,x756 } )+$signed( -{ 2'b0,x245 }<<<3'd1 )+$signed( { 3'b0,x501 }<<<3'd2 )+$signed( -{ 2'b0,x757 }<<<3'd1 )+$signed(11'd32);
assign y314=temp_y[314][11] ==1'b1 ? 5'd0 :  
        temp_y[314][8] ==1'b1 ? 5'd31 : 
        temp_y[314][2]==1'b1 ? temp_y[314][7:3]+1'b1 : temp_y[314][7:3];
assign temp_y[378] = 
+$signed( -{ 1'b0,x228 } )+$signed( -{ 2'b0,x484 }<<<3'd1 )+$signed( -{ 1'b0,x740 } )+$signed( { 1'b0,x229 }  )+$signed( { 2'b0,x485 } <<<3'd1 )+$signed( { 1'b0,x741 }  )+$signed( { 1'b0,x244 }  )+$signed( { 2'b0,x500 } <<<3'd1 )+$signed( { 2'b0,x756 } <<<3'd1 )+$signed( -{ 1'b0,x245 } )+$signed( -{ 2'b0,x501 }<<<3'd1 )+$signed( -{ 1'b0,x757 } )-$signed(11'd68);
assign y378=temp_y[378][11] ==1'b1 ? 5'd0 :  
        temp_y[378][8] ==1'b1 ? 5'd31 : 
        temp_y[378][2]==1'b1 ? temp_y[378][7:3]+1'b1 : temp_y[378][7:3];
assign temp_y[442] = 
+$signed( { 1'b0,x484 }  )+$signed( { 1'b0,x741 }  )+$signed( { 1'b0,x757 }  )-$signed(11'd108);
assign y442=temp_y[442][11] ==1'b1 ? 5'd0 :  
        temp_y[442][8] ==1'b1 ? 5'd31 : 
        temp_y[442][2]==1'b1 ? temp_y[442][7:3]+1'b1 : temp_y[442][7:3];
assign temp_y[506] = 
+$signed( -{ 2'b0,x228 }<<<3'd1 )+$signed( { 2'b0,x740 } <<<3'd1 )+$signed( -{ 2'b0,x229 }<<<3'd1 )+$signed( { 1'b0,x485 }  )+$signed( { 1'b0,x741 }  )+$signed( -{ 2'b0,x244 }<<<3'd1 )+$signed( { 1'b0,x500 }  )+$signed( { 1'b0,x756 }  )+$signed( -{ 1'b0,x245 } )+$signed(11'd64);
assign y506=temp_y[506][11] ==1'b1 ? 5'd0 :  
        temp_y[506][8] ==1'b1 ? 5'd31 : 
        temp_y[506][2]==1'b1 ? temp_y[506][7:3]+1'b1 : temp_y[506][7:3];
assign temp_y[570] = 
+$signed( -{ 2'b0,x228 }<<<3'd1 )+$signed( -{ 1'b0,x484 } )+$signed( -{ 3'b0,x229 }<<<3'd2)+$signed( { 1'b0,x244 }  )+$signed( { 1'b0,x500 }  )+$signed( { 3'b0,x245 }<<<3'd2 )+$signed(11'd16);
assign y570=temp_y[570][11] ==1'b1 ? 5'd0 :  
        temp_y[570][8] ==1'b1 ? 5'd31 : 
        temp_y[570][2]==1'b1 ? temp_y[570][7:3]+1'b1 : temp_y[570][7:3];
assign temp_y[634] = 
+$signed( { 2'b0,x484 } <<<3'd1 )+$signed( { 2'b0,x740 } <<<3'd1 )+$signed( -{ 1'b0,x229 } )+$signed( -{ 2'b0,x485 }<<<3'd1 )+$signed( -{ 2'b0,x741 }<<<3'd1 )+$signed( { 2'b0,x500 } <<<3'd1 )+$signed( { 1'b0,x756 }  )+$signed( -{ 2'b0,x501 }<<<3'd1 )-$signed(11'd8);
assign y634=temp_y[634][11] ==1'b1 ? 5'd0 :  
        temp_y[634][8] ==1'b1 ? 5'd31 : 
        temp_y[634][2]==1'b1 ? temp_y[634][7:3]+1'b1 : temp_y[634][7:3];
assign temp_y[59] = 
+$signed( -{ 2'b0,x486 }<<<3'd1 )+$signed( -{ 1'b0,x742 } )+$signed( { 1'b0,x231 }  )+$signed( { 1'b0,x487 }  )+$signed( { 1'b0,x743 }  )+$signed( -{ 2'b0,x502 }<<<3'd1 )+$signed( -{ 2'b0,x758 }<<<3'd1 )+$signed( { 2'b0,x503 } <<<3'd1 )+$signed( { 2'b0,x759 } <<<3'd1 )-$signed(11'd16);
assign y59=temp_y[59][11] ==1'b1 ? 5'd0 :  
        temp_y[59][8] ==1'b1 ? 5'd31 : 
        temp_y[59][2]==1'b1 ? temp_y[59][7:3]+1'b1 : temp_y[59][7:3];
assign temp_y[123] = 
+$signed( { 3'b0,x230 }<<<3'd2 )+$signed( -{ 2'b0,x486 }<<<3'd1 )+$signed( -{ 2'b0,x742 }<<<3'd1 )+$signed( { 2'b0,x231 } <<<3'd1 )+$signed( -{ 3'b0,x487 }<<<3'd2)+$signed( { 1'b0,x743 }  )+$signed( -{ 1'b0,x246 } )+$signed( { 1'b0,x758 }  )+$signed( -{ 2'b0,x247 }<<<3'd1 )+$signed( -{ 1'b0,x503 } )+$signed( { 2'b0,x759 } <<<3'd1 )+$signed(11'd24);
assign y123=temp_y[123][11] ==1'b1 ? 5'd0 :  
        temp_y[123][8] ==1'b1 ? 5'd31 : 
        temp_y[123][2]==1'b1 ? temp_y[123][7:3]+1'b1 : temp_y[123][7:3];
assign temp_y[187] = 
+$signed( { 2'b0,x230 } <<<3'd1 )+$signed( { 2'b0,x486 } <<<3'd1 )+$signed( { 1'b0,x742 }  )+$signed( { 2'b0,x231 } <<<3'd1 )+$signed( -{ 1'b0,x487 } )+$signed( { 1'b0,x743 }  )+$signed( -{ 2'b0,x246 }<<<3'd1 )+$signed( -{ 2'b0,x502 }<<<3'd1 )+$signed( -{ 1'b0,x758 } )+$signed( -{ 1'b0,x247 } )+$signed( -{ 1'b0,x503 } )+$signed( -{ 1'b0,x759 } )+$signed(11'd16);
assign y187=temp_y[187][11] ==1'b1 ? 5'd0 :  
        temp_y[187][8] ==1'b1 ? 5'd31 : 
        temp_y[187][2]==1'b1 ? temp_y[187][7:3]+1'b1 : temp_y[187][7:3];
assign temp_y[251] = 
+$signed( { 1'b0,x230 }  )+$signed( -{ 1'b0,x486 } )+$signed( { 1'b0,x231 }  )+$signed( -{ 1'b0,x487 } )+$signed( { 2'b0,x246 } <<<3'd1 )+$signed( -{ 1'b0,x502 } )+$signed( -{ 1'b0,x758 } )+$signed( { 2'b0,x247 } <<<3'd1 )+$signed( -{ 1'b0,x503 } )+$signed( -{ 2'b0,x759 }<<<3'd1 )+$signed(11'd40);
assign y251=temp_y[251][11] ==1'b1 ? 5'd0 :  
        temp_y[251][8] ==1'b1 ? 5'd31 : 
        temp_y[251][2]==1'b1 ? temp_y[251][7:3]+1'b1 : temp_y[251][7:3];
assign temp_y[315] = 
+$signed( -{ 1'b0,x230 } )+$signed( { 2'b0,x486 } <<<3'd1 )+$signed( -{ 1'b0,x742 } )+$signed( -{ 1'b0,x231 } )+$signed( { 2'b0,x487 } <<<3'd1 )+$signed( -{ 2'b0,x743 }<<<3'd1 )+$signed( -{ 1'b0,x246 } )+$signed( { 2'b0,x502 } <<<3'd1 )+$signed( -{ 1'b0,x758 } )+$signed( -{ 2'b0,x247 }<<<3'd1 )+$signed( { 3'b0,x503 }<<<3'd2 )+$signed( -{ 2'b0,x759 }<<<3'd1 )+$signed(11'd32);
assign y315=temp_y[315][11] ==1'b1 ? 5'd0 :  
        temp_y[315][8] ==1'b1 ? 5'd31 : 
        temp_y[315][2]==1'b1 ? temp_y[315][7:3]+1'b1 : temp_y[315][7:3];
assign temp_y[379] = 
+$signed( -{ 1'b0,x230 } )+$signed( -{ 2'b0,x486 }<<<3'd1 )+$signed( -{ 1'b0,x742 } )+$signed( { 1'b0,x231 }  )+$signed( { 2'b0,x487 } <<<3'd1 )+$signed( { 1'b0,x743 }  )+$signed( { 1'b0,x246 }  )+$signed( { 2'b0,x502 } <<<3'd1 )+$signed( { 2'b0,x758 } <<<3'd1 )+$signed( -{ 1'b0,x247 } )+$signed( -{ 2'b0,x503 }<<<3'd1 )+$signed( -{ 1'b0,x759 } )-$signed(11'd68);
assign y379=temp_y[379][11] ==1'b1 ? 5'd0 :  
        temp_y[379][8] ==1'b1 ? 5'd31 : 
        temp_y[379][2]==1'b1 ? temp_y[379][7:3]+1'b1 : temp_y[379][7:3];
assign temp_y[443] = 
+$signed( { 1'b0,x486 }  )+$signed( { 1'b0,x743 }  )+$signed( { 1'b0,x759 }  )-$signed(11'd108);
assign y443=temp_y[443][11] ==1'b1 ? 5'd0 :  
        temp_y[443][8] ==1'b1 ? 5'd31 : 
        temp_y[443][2]==1'b1 ? temp_y[443][7:3]+1'b1 : temp_y[443][7:3];
assign temp_y[507] = 
+$signed( -{ 2'b0,x230 }<<<3'd1 )+$signed( { 2'b0,x742 } <<<3'd1 )+$signed( -{ 2'b0,x231 }<<<3'd1 )+$signed( { 1'b0,x487 }  )+$signed( { 1'b0,x743 }  )+$signed( -{ 2'b0,x246 }<<<3'd1 )+$signed( { 1'b0,x502 }  )+$signed( { 1'b0,x758 }  )+$signed( -{ 1'b0,x247 } )+$signed(11'd64);
assign y507=temp_y[507][11] ==1'b1 ? 5'd0 :  
        temp_y[507][8] ==1'b1 ? 5'd31 : 
        temp_y[507][2]==1'b1 ? temp_y[507][7:3]+1'b1 : temp_y[507][7:3];
assign temp_y[571] = 
+$signed( -{ 2'b0,x230 }<<<3'd1 )+$signed( -{ 1'b0,x486 } )+$signed( -{ 3'b0,x231 }<<<3'd2)+$signed( { 1'b0,x246 }  )+$signed( { 1'b0,x502 }  )+$signed( { 3'b0,x247 }<<<3'd2 )+$signed(11'd16);
assign y571=temp_y[571][11] ==1'b1 ? 5'd0 :  
        temp_y[571][8] ==1'b1 ? 5'd31 : 
        temp_y[571][2]==1'b1 ? temp_y[571][7:3]+1'b1 : temp_y[571][7:3];
assign temp_y[635] = 
+$signed( { 2'b0,x486 } <<<3'd1 )+$signed( { 2'b0,x742 } <<<3'd1 )+$signed( -{ 1'b0,x231 } )+$signed( -{ 2'b0,x487 }<<<3'd1 )+$signed( -{ 2'b0,x743 }<<<3'd1 )+$signed( { 2'b0,x502 } <<<3'd1 )+$signed( { 1'b0,x758 }  )+$signed( -{ 2'b0,x503 }<<<3'd1 )-$signed(11'd8);
assign y635=temp_y[635][11] ==1'b1 ? 5'd0 :  
        temp_y[635][8] ==1'b1 ? 5'd31 : 
        temp_y[635][2]==1'b1 ? temp_y[635][7:3]+1'b1 : temp_y[635][7:3];
assign temp_y[60] = 
+$signed( -{ 2'b0,x488 }<<<3'd1 )+$signed( -{ 1'b0,x744 } )+$signed( { 1'b0,x233 }  )+$signed( { 1'b0,x489 }  )+$signed( { 1'b0,x745 }  )+$signed( -{ 2'b0,x504 }<<<3'd1 )+$signed( -{ 2'b0,x760 }<<<3'd1 )+$signed( { 2'b0,x505 } <<<3'd1 )+$signed( { 2'b0,x761 } <<<3'd1 )-$signed(11'd16);
assign y60=temp_y[60][11] ==1'b1 ? 5'd0 :  
        temp_y[60][8] ==1'b1 ? 5'd31 : 
        temp_y[60][2]==1'b1 ? temp_y[60][7:3]+1'b1 : temp_y[60][7:3];
assign temp_y[124] = 
+$signed( { 3'b0,x232 }<<<3'd2 )+$signed( -{ 2'b0,x488 }<<<3'd1 )+$signed( -{ 2'b0,x744 }<<<3'd1 )+$signed( { 2'b0,x233 } <<<3'd1 )+$signed( -{ 3'b0,x489 }<<<3'd2)+$signed( { 1'b0,x745 }  )+$signed( -{ 1'b0,x248 } )+$signed( { 1'b0,x760 }  )+$signed( -{ 2'b0,x249 }<<<3'd1 )+$signed( -{ 1'b0,x505 } )+$signed( { 2'b0,x761 } <<<3'd1 )+$signed(11'd24);
assign y124=temp_y[124][11] ==1'b1 ? 5'd0 :  
        temp_y[124][8] ==1'b1 ? 5'd31 : 
        temp_y[124][2]==1'b1 ? temp_y[124][7:3]+1'b1 : temp_y[124][7:3];
assign temp_y[188] = 
+$signed( { 2'b0,x232 } <<<3'd1 )+$signed( { 2'b0,x488 } <<<3'd1 )+$signed( { 1'b0,x744 }  )+$signed( { 2'b0,x233 } <<<3'd1 )+$signed( -{ 1'b0,x489 } )+$signed( { 1'b0,x745 }  )+$signed( -{ 2'b0,x248 }<<<3'd1 )+$signed( -{ 2'b0,x504 }<<<3'd1 )+$signed( -{ 1'b0,x760 } )+$signed( -{ 1'b0,x249 } )+$signed( -{ 1'b0,x505 } )+$signed( -{ 1'b0,x761 } )+$signed(11'd16);
assign y188=temp_y[188][11] ==1'b1 ? 5'd0 :  
        temp_y[188][8] ==1'b1 ? 5'd31 : 
        temp_y[188][2]==1'b1 ? temp_y[188][7:3]+1'b1 : temp_y[188][7:3];
assign temp_y[252] = 
+$signed( { 1'b0,x232 }  )+$signed( -{ 1'b0,x488 } )+$signed( { 1'b0,x233 }  )+$signed( -{ 1'b0,x489 } )+$signed( { 2'b0,x248 } <<<3'd1 )+$signed( -{ 1'b0,x504 } )+$signed( -{ 1'b0,x760 } )+$signed( { 2'b0,x249 } <<<3'd1 )+$signed( -{ 1'b0,x505 } )+$signed( -{ 2'b0,x761 }<<<3'd1 )+$signed(11'd40);
assign y252=temp_y[252][11] ==1'b1 ? 5'd0 :  
        temp_y[252][8] ==1'b1 ? 5'd31 : 
        temp_y[252][2]==1'b1 ? temp_y[252][7:3]+1'b1 : temp_y[252][7:3];
assign temp_y[316] = 
+$signed( -{ 1'b0,x232 } )+$signed( { 2'b0,x488 } <<<3'd1 )+$signed( -{ 1'b0,x744 } )+$signed( -{ 1'b0,x233 } )+$signed( { 2'b0,x489 } <<<3'd1 )+$signed( -{ 2'b0,x745 }<<<3'd1 )+$signed( -{ 1'b0,x248 } )+$signed( { 2'b0,x504 } <<<3'd1 )+$signed( -{ 1'b0,x760 } )+$signed( -{ 2'b0,x249 }<<<3'd1 )+$signed( { 3'b0,x505 }<<<3'd2 )+$signed( -{ 2'b0,x761 }<<<3'd1 )+$signed(11'd32);
assign y316=temp_y[316][11] ==1'b1 ? 5'd0 :  
        temp_y[316][8] ==1'b1 ? 5'd31 : 
        temp_y[316][2]==1'b1 ? temp_y[316][7:3]+1'b1 : temp_y[316][7:3];
assign temp_y[380] = 
+$signed( -{ 1'b0,x232 } )+$signed( -{ 2'b0,x488 }<<<3'd1 )+$signed( -{ 1'b0,x744 } )+$signed( { 1'b0,x233 }  )+$signed( { 2'b0,x489 } <<<3'd1 )+$signed( { 1'b0,x745 }  )+$signed( { 1'b0,x248 }  )+$signed( { 2'b0,x504 } <<<3'd1 )+$signed( { 2'b0,x760 } <<<3'd1 )+$signed( -{ 1'b0,x249 } )+$signed( -{ 2'b0,x505 }<<<3'd1 )+$signed( -{ 1'b0,x761 } )-$signed(11'd68);
assign y380=temp_y[380][11] ==1'b1 ? 5'd0 :  
        temp_y[380][8] ==1'b1 ? 5'd31 : 
        temp_y[380][2]==1'b1 ? temp_y[380][7:3]+1'b1 : temp_y[380][7:3];
assign temp_y[444] = 
+$signed( { 1'b0,x488 }  )+$signed( { 1'b0,x745 }  )+$signed( { 1'b0,x761 }  )-$signed(11'd108);
assign y444=temp_y[444][11] ==1'b1 ? 5'd0 :  
        temp_y[444][8] ==1'b1 ? 5'd31 : 
        temp_y[444][2]==1'b1 ? temp_y[444][7:3]+1'b1 : temp_y[444][7:3];
assign temp_y[508] = 
+$signed( -{ 2'b0,x232 }<<<3'd1 )+$signed( { 2'b0,x744 } <<<3'd1 )+$signed( -{ 2'b0,x233 }<<<3'd1 )+$signed( { 1'b0,x489 }  )+$signed( { 1'b0,x745 }  )+$signed( -{ 2'b0,x248 }<<<3'd1 )+$signed( { 1'b0,x504 }  )+$signed( { 1'b0,x760 }  )+$signed( -{ 1'b0,x249 } )+$signed(11'd64);
assign y508=temp_y[508][11] ==1'b1 ? 5'd0 :  
        temp_y[508][8] ==1'b1 ? 5'd31 : 
        temp_y[508][2]==1'b1 ? temp_y[508][7:3]+1'b1 : temp_y[508][7:3];
assign temp_y[572] = 
+$signed( -{ 2'b0,x232 }<<<3'd1 )+$signed( -{ 1'b0,x488 } )+$signed( -{ 3'b0,x233 }<<<3'd2)+$signed( { 1'b0,x248 }  )+$signed( { 1'b0,x504 }  )+$signed( { 3'b0,x249 }<<<3'd2 )+$signed(11'd16);
assign y572=temp_y[572][11] ==1'b1 ? 5'd0 :  
        temp_y[572][8] ==1'b1 ? 5'd31 : 
        temp_y[572][2]==1'b1 ? temp_y[572][7:3]+1'b1 : temp_y[572][7:3];
assign temp_y[636] = 
+$signed( { 2'b0,x488 } <<<3'd1 )+$signed( { 2'b0,x744 } <<<3'd1 )+$signed( -{ 1'b0,x233 } )+$signed( -{ 2'b0,x489 }<<<3'd1 )+$signed( -{ 2'b0,x745 }<<<3'd1 )+$signed( { 2'b0,x504 } <<<3'd1 )+$signed( { 1'b0,x760 }  )+$signed( -{ 2'b0,x505 }<<<3'd1 )-$signed(11'd8);
assign y636=temp_y[636][11] ==1'b1 ? 5'd0 :  
        temp_y[636][8] ==1'b1 ? 5'd31 : 
        temp_y[636][2]==1'b1 ? temp_y[636][7:3]+1'b1 : temp_y[636][7:3];
assign temp_y[61] = 
+$signed( -{ 2'b0,x490 }<<<3'd1 )+$signed( -{ 1'b0,x746 } )+$signed( { 1'b0,x235 }  )+$signed( { 1'b0,x491 }  )+$signed( { 1'b0,x747 }  )+$signed( -{ 2'b0,x506 }<<<3'd1 )+$signed( -{ 2'b0,x762 }<<<3'd1 )+$signed( { 2'b0,x507 } <<<3'd1 )+$signed( { 2'b0,x763 } <<<3'd1 )-$signed(11'd16);
assign y61=temp_y[61][11] ==1'b1 ? 5'd0 :  
        temp_y[61][8] ==1'b1 ? 5'd31 : 
        temp_y[61][2]==1'b1 ? temp_y[61][7:3]+1'b1 : temp_y[61][7:3];
assign temp_y[125] = 
+$signed( { 3'b0,x234 }<<<3'd2 )+$signed( -{ 2'b0,x490 }<<<3'd1 )+$signed( -{ 2'b0,x746 }<<<3'd1 )+$signed( { 2'b0,x235 } <<<3'd1 )+$signed( -{ 3'b0,x491 }<<<3'd2)+$signed( { 1'b0,x747 }  )+$signed( -{ 1'b0,x250 } )+$signed( { 1'b0,x762 }  )+$signed( -{ 2'b0,x251 }<<<3'd1 )+$signed( -{ 1'b0,x507 } )+$signed( { 2'b0,x763 } <<<3'd1 )+$signed(11'd24);
assign y125=temp_y[125][11] ==1'b1 ? 5'd0 :  
        temp_y[125][8] ==1'b1 ? 5'd31 : 
        temp_y[125][2]==1'b1 ? temp_y[125][7:3]+1'b1 : temp_y[125][7:3];
assign temp_y[189] = 
+$signed( { 2'b0,x234 } <<<3'd1 )+$signed( { 2'b0,x490 } <<<3'd1 )+$signed( { 1'b0,x746 }  )+$signed( { 2'b0,x235 } <<<3'd1 )+$signed( -{ 1'b0,x491 } )+$signed( { 1'b0,x747 }  )+$signed( -{ 2'b0,x250 }<<<3'd1 )+$signed( -{ 2'b0,x506 }<<<3'd1 )+$signed( -{ 1'b0,x762 } )+$signed( -{ 1'b0,x251 } )+$signed( -{ 1'b0,x507 } )+$signed( -{ 1'b0,x763 } )+$signed(11'd16);
assign y189=temp_y[189][11] ==1'b1 ? 5'd0 :  
        temp_y[189][8] ==1'b1 ? 5'd31 : 
        temp_y[189][2]==1'b1 ? temp_y[189][7:3]+1'b1 : temp_y[189][7:3];
assign temp_y[253] = 
+$signed( { 1'b0,x234 }  )+$signed( -{ 1'b0,x490 } )+$signed( { 1'b0,x235 }  )+$signed( -{ 1'b0,x491 } )+$signed( { 2'b0,x250 } <<<3'd1 )+$signed( -{ 1'b0,x506 } )+$signed( -{ 1'b0,x762 } )+$signed( { 2'b0,x251 } <<<3'd1 )+$signed( -{ 1'b0,x507 } )+$signed( -{ 2'b0,x763 }<<<3'd1 )+$signed(11'd40);
assign y253=temp_y[253][11] ==1'b1 ? 5'd0 :  
        temp_y[253][8] ==1'b1 ? 5'd31 : 
        temp_y[253][2]==1'b1 ? temp_y[253][7:3]+1'b1 : temp_y[253][7:3];
assign temp_y[317] = 
+$signed( -{ 1'b0,x234 } )+$signed( { 2'b0,x490 } <<<3'd1 )+$signed( -{ 1'b0,x746 } )+$signed( -{ 1'b0,x235 } )+$signed( { 2'b0,x491 } <<<3'd1 )+$signed( -{ 2'b0,x747 }<<<3'd1 )+$signed( -{ 1'b0,x250 } )+$signed( { 2'b0,x506 } <<<3'd1 )+$signed( -{ 1'b0,x762 } )+$signed( -{ 2'b0,x251 }<<<3'd1 )+$signed( { 3'b0,x507 }<<<3'd2 )+$signed( -{ 2'b0,x763 }<<<3'd1 )+$signed(11'd32);
assign y317=temp_y[317][11] ==1'b1 ? 5'd0 :  
        temp_y[317][8] ==1'b1 ? 5'd31 : 
        temp_y[317][2]==1'b1 ? temp_y[317][7:3]+1'b1 : temp_y[317][7:3];
assign temp_y[381] = 
+$signed( -{ 1'b0,x234 } )+$signed( -{ 2'b0,x490 }<<<3'd1 )+$signed( -{ 1'b0,x746 } )+$signed( { 1'b0,x235 }  )+$signed( { 2'b0,x491 } <<<3'd1 )+$signed( { 1'b0,x747 }  )+$signed( { 1'b0,x250 }  )+$signed( { 2'b0,x506 } <<<3'd1 )+$signed( { 2'b0,x762 } <<<3'd1 )+$signed( -{ 1'b0,x251 } )+$signed( -{ 2'b0,x507 }<<<3'd1 )+$signed( -{ 1'b0,x763 } )-$signed(11'd68);
assign y381=temp_y[381][11] ==1'b1 ? 5'd0 :  
        temp_y[381][8] ==1'b1 ? 5'd31 : 
        temp_y[381][2]==1'b1 ? temp_y[381][7:3]+1'b1 : temp_y[381][7:3];
assign temp_y[445] = 
+$signed( { 1'b0,x490 }  )+$signed( { 1'b0,x747 }  )+$signed( { 1'b0,x763 }  )-$signed(11'd108);
assign y445=temp_y[445][11] ==1'b1 ? 5'd0 :  
        temp_y[445][8] ==1'b1 ? 5'd31 : 
        temp_y[445][2]==1'b1 ? temp_y[445][7:3]+1'b1 : temp_y[445][7:3];
assign temp_y[509] = 
+$signed( -{ 2'b0,x234 }<<<3'd1 )+$signed( { 2'b0,x746 } <<<3'd1 )+$signed( -{ 2'b0,x235 }<<<3'd1 )+$signed( { 1'b0,x491 }  )+$signed( { 1'b0,x747 }  )+$signed( -{ 2'b0,x250 }<<<3'd1 )+$signed( { 1'b0,x506 }  )+$signed( { 1'b0,x762 }  )+$signed( -{ 1'b0,x251 } )+$signed(11'd64);
assign y509=temp_y[509][11] ==1'b1 ? 5'd0 :  
        temp_y[509][8] ==1'b1 ? 5'd31 : 
        temp_y[509][2]==1'b1 ? temp_y[509][7:3]+1'b1 : temp_y[509][7:3];
assign temp_y[573] = 
+$signed( -{ 2'b0,x234 }<<<3'd1 )+$signed( -{ 1'b0,x490 } )+$signed( -{ 3'b0,x235 }<<<3'd2)+$signed( { 1'b0,x250 }  )+$signed( { 1'b0,x506 }  )+$signed( { 3'b0,x251 }<<<3'd2 )+$signed(11'd16);
assign y573=temp_y[573][11] ==1'b1 ? 5'd0 :  
        temp_y[573][8] ==1'b1 ? 5'd31 : 
        temp_y[573][2]==1'b1 ? temp_y[573][7:3]+1'b1 : temp_y[573][7:3];
assign temp_y[637] = 
+$signed( { 2'b0,x490 } <<<3'd1 )+$signed( { 2'b0,x746 } <<<3'd1 )+$signed( -{ 1'b0,x235 } )+$signed( -{ 2'b0,x491 }<<<3'd1 )+$signed( -{ 2'b0,x747 }<<<3'd1 )+$signed( { 2'b0,x506 } <<<3'd1 )+$signed( { 1'b0,x762 }  )+$signed( -{ 2'b0,x507 }<<<3'd1 )-$signed(11'd8);
assign y637=temp_y[637][11] ==1'b1 ? 5'd0 :  
        temp_y[637][8] ==1'b1 ? 5'd31 : 
        temp_y[637][2]==1'b1 ? temp_y[637][7:3]+1'b1 : temp_y[637][7:3];
assign temp_y[62] = 
+$signed( -{ 2'b0,x492 }<<<3'd1 )+$signed( -{ 1'b0,x748 } )+$signed( { 1'b0,x237 }  )+$signed( { 1'b0,x493 }  )+$signed( { 1'b0,x749 }  )+$signed( -{ 2'b0,x508 }<<<3'd1 )+$signed( -{ 2'b0,x764 }<<<3'd1 )+$signed( { 2'b0,x509 } <<<3'd1 )+$signed( { 2'b0,x765 } <<<3'd1 )-$signed(11'd16);
assign y62=temp_y[62][11] ==1'b1 ? 5'd0 :  
        temp_y[62][8] ==1'b1 ? 5'd31 : 
        temp_y[62][2]==1'b1 ? temp_y[62][7:3]+1'b1 : temp_y[62][7:3];
assign temp_y[126] = 
+$signed( { 3'b0,x236 }<<<3'd2 )+$signed( -{ 2'b0,x492 }<<<3'd1 )+$signed( -{ 2'b0,x748 }<<<3'd1 )+$signed( { 2'b0,x237 } <<<3'd1 )+$signed( -{ 3'b0,x493 }<<<3'd2)+$signed( { 1'b0,x749 }  )+$signed( -{ 1'b0,x252 } )+$signed( { 1'b0,x764 }  )+$signed( -{ 2'b0,x253 }<<<3'd1 )+$signed( -{ 1'b0,x509 } )+$signed( { 2'b0,x765 } <<<3'd1 )+$signed(11'd24);
assign y126=temp_y[126][11] ==1'b1 ? 5'd0 :  
        temp_y[126][8] ==1'b1 ? 5'd31 : 
        temp_y[126][2]==1'b1 ? temp_y[126][7:3]+1'b1 : temp_y[126][7:3];
assign temp_y[190] = 
+$signed( { 2'b0,x236 } <<<3'd1 )+$signed( { 2'b0,x492 } <<<3'd1 )+$signed( { 1'b0,x748 }  )+$signed( { 2'b0,x237 } <<<3'd1 )+$signed( -{ 1'b0,x493 } )+$signed( { 1'b0,x749 }  )+$signed( -{ 2'b0,x252 }<<<3'd1 )+$signed( -{ 2'b0,x508 }<<<3'd1 )+$signed( -{ 1'b0,x764 } )+$signed( -{ 1'b0,x253 } )+$signed( -{ 1'b0,x509 } )+$signed( -{ 1'b0,x765 } )+$signed(11'd16);
assign y190=temp_y[190][11] ==1'b1 ? 5'd0 :  
        temp_y[190][8] ==1'b1 ? 5'd31 : 
        temp_y[190][2]==1'b1 ? temp_y[190][7:3]+1'b1 : temp_y[190][7:3];
assign temp_y[254] = 
+$signed( { 1'b0,x236 }  )+$signed( -{ 1'b0,x492 } )+$signed( { 1'b0,x237 }  )+$signed( -{ 1'b0,x493 } )+$signed( { 2'b0,x252 } <<<3'd1 )+$signed( -{ 1'b0,x508 } )+$signed( -{ 1'b0,x764 } )+$signed( { 2'b0,x253 } <<<3'd1 )+$signed( -{ 1'b0,x509 } )+$signed( -{ 2'b0,x765 }<<<3'd1 )+$signed(11'd40);
assign y254=temp_y[254][11] ==1'b1 ? 5'd0 :  
        temp_y[254][8] ==1'b1 ? 5'd31 : 
        temp_y[254][2]==1'b1 ? temp_y[254][7:3]+1'b1 : temp_y[254][7:3];
assign temp_y[318] = 
+$signed( -{ 1'b0,x236 } )+$signed( { 2'b0,x492 } <<<3'd1 )+$signed( -{ 1'b0,x748 } )+$signed( -{ 1'b0,x237 } )+$signed( { 2'b0,x493 } <<<3'd1 )+$signed( -{ 2'b0,x749 }<<<3'd1 )+$signed( -{ 1'b0,x252 } )+$signed( { 2'b0,x508 } <<<3'd1 )+$signed( -{ 1'b0,x764 } )+$signed( -{ 2'b0,x253 }<<<3'd1 )+$signed( { 3'b0,x509 }<<<3'd2 )+$signed( -{ 2'b0,x765 }<<<3'd1 )+$signed(11'd32);
assign y318=temp_y[318][11] ==1'b1 ? 5'd0 :  
        temp_y[318][8] ==1'b1 ? 5'd31 : 
        temp_y[318][2]==1'b1 ? temp_y[318][7:3]+1'b1 : temp_y[318][7:3];
assign temp_y[382] = 
+$signed( -{ 1'b0,x236 } )+$signed( -{ 2'b0,x492 }<<<3'd1 )+$signed( -{ 1'b0,x748 } )+$signed( { 1'b0,x237 }  )+$signed( { 2'b0,x493 } <<<3'd1 )+$signed( { 1'b0,x749 }  )+$signed( { 1'b0,x252 }  )+$signed( { 2'b0,x508 } <<<3'd1 )+$signed( { 2'b0,x764 } <<<3'd1 )+$signed( -{ 1'b0,x253 } )+$signed( -{ 2'b0,x509 }<<<3'd1 )+$signed( -{ 1'b0,x765 } )-$signed(11'd68);
assign y382=temp_y[382][11] ==1'b1 ? 5'd0 :  
        temp_y[382][8] ==1'b1 ? 5'd31 : 
        temp_y[382][2]==1'b1 ? temp_y[382][7:3]+1'b1 : temp_y[382][7:3];
assign temp_y[446] = 
+$signed( { 1'b0,x492 }  )+$signed( { 1'b0,x749 }  )+$signed( { 1'b0,x765 }  )-$signed(11'd108);
assign y446=temp_y[446][11] ==1'b1 ? 5'd0 :  
        temp_y[446][8] ==1'b1 ? 5'd31 : 
        temp_y[446][2]==1'b1 ? temp_y[446][7:3]+1'b1 : temp_y[446][7:3];
assign temp_y[510] = 
+$signed( -{ 2'b0,x236 }<<<3'd1 )+$signed( { 2'b0,x748 } <<<3'd1 )+$signed( -{ 2'b0,x237 }<<<3'd1 )+$signed( { 1'b0,x493 }  )+$signed( { 1'b0,x749 }  )+$signed( -{ 2'b0,x252 }<<<3'd1 )+$signed( { 1'b0,x508 }  )+$signed( { 1'b0,x764 }  )+$signed( -{ 1'b0,x253 } )+$signed(11'd64);
assign y510=temp_y[510][11] ==1'b1 ? 5'd0 :  
        temp_y[510][8] ==1'b1 ? 5'd31 : 
        temp_y[510][2]==1'b1 ? temp_y[510][7:3]+1'b1 : temp_y[510][7:3];
assign temp_y[574] = 
+$signed( -{ 2'b0,x236 }<<<3'd1 )+$signed( -{ 1'b0,x492 } )+$signed( -{ 3'b0,x237 }<<<3'd2)+$signed( { 1'b0,x252 }  )+$signed( { 1'b0,x508 }  )+$signed( { 3'b0,x253 }<<<3'd2 )+$signed(11'd16);
assign y574=temp_y[574][11] ==1'b1 ? 5'd0 :  
        temp_y[574][8] ==1'b1 ? 5'd31 : 
        temp_y[574][2]==1'b1 ? temp_y[574][7:3]+1'b1 : temp_y[574][7:3];
assign temp_y[638] = 
+$signed( { 2'b0,x492 } <<<3'd1 )+$signed( { 2'b0,x748 } <<<3'd1 )+$signed( -{ 1'b0,x237 } )+$signed( -{ 2'b0,x493 }<<<3'd1 )+$signed( -{ 2'b0,x749 }<<<3'd1 )+$signed( { 2'b0,x508 } <<<3'd1 )+$signed( { 1'b0,x764 }  )+$signed( -{ 2'b0,x509 }<<<3'd1 )-$signed(11'd8);
assign y638=temp_y[638][11] ==1'b1 ? 5'd0 :  
        temp_y[638][8] ==1'b1 ? 5'd31 : 
        temp_y[638][2]==1'b1 ? temp_y[638][7:3]+1'b1 : temp_y[638][7:3];
assign temp_y[63] = 
+$signed( -{ 2'b0,x494 }<<<3'd1 )+$signed( -{ 1'b0,x750 } )+$signed( { 1'b0,x239 }  )+$signed( { 1'b0,x495 }  )+$signed( { 1'b0,x751 }  )+$signed( -{ 2'b0,x510 }<<<3'd1 )+$signed( -{ 2'b0,x766 }<<<3'd1 )+$signed( { 2'b0,x511 } <<<3'd1 )+$signed( { 2'b0,x767 } <<<3'd1 )-$signed(11'd16);
assign y63=temp_y[63][11] ==1'b1 ? 5'd0 :  
        temp_y[63][8] ==1'b1 ? 5'd31 : 
        temp_y[63][2]==1'b1 ? temp_y[63][7:3]+1'b1 : temp_y[63][7:3];
assign temp_y[127] = 
+$signed( { 3'b0,x238 }<<<3'd2 )+$signed( -{ 2'b0,x494 }<<<3'd1 )+$signed( -{ 2'b0,x750 }<<<3'd1 )+$signed( { 2'b0,x239 } <<<3'd1 )+$signed( -{ 3'b0,x495 }<<<3'd2)+$signed( { 1'b0,x751 }  )+$signed( -{ 1'b0,x254 } )+$signed( { 1'b0,x766 }  )+$signed( -{ 2'b0,x255 }<<<3'd1 )+$signed( -{ 1'b0,x511 } )+$signed( { 2'b0,x767 } <<<3'd1 )+$signed(11'd24);
assign y127=temp_y[127][11] ==1'b1 ? 5'd0 :  
        temp_y[127][8] ==1'b1 ? 5'd31 : 
        temp_y[127][2]==1'b1 ? temp_y[127][7:3]+1'b1 : temp_y[127][7:3];
assign temp_y[191] = 
+$signed( { 2'b0,x238 } <<<3'd1 )+$signed( { 2'b0,x494 } <<<3'd1 )+$signed( { 1'b0,x750 }  )+$signed( { 2'b0,x239 } <<<3'd1 )+$signed( -{ 1'b0,x495 } )+$signed( { 1'b0,x751 }  )+$signed( -{ 2'b0,x254 }<<<3'd1 )+$signed( -{ 2'b0,x510 }<<<3'd1 )+$signed( -{ 1'b0,x766 } )+$signed( -{ 1'b0,x255 } )+$signed( -{ 1'b0,x511 } )+$signed( -{ 1'b0,x767 } )+$signed(11'd16);
assign y191=temp_y[191][11] ==1'b1 ? 5'd0 :  
        temp_y[191][8] ==1'b1 ? 5'd31 : 
        temp_y[191][2]==1'b1 ? temp_y[191][7:3]+1'b1 : temp_y[191][7:3];
assign temp_y[255] = 
+$signed( { 1'b0,x238 }  )+$signed( -{ 1'b0,x494 } )+$signed( { 1'b0,x239 }  )+$signed( -{ 1'b0,x495 } )+$signed( { 2'b0,x254 } <<<3'd1 )+$signed( -{ 1'b0,x510 } )+$signed( -{ 1'b0,x766 } )+$signed( { 2'b0,x255 } <<<3'd1 )+$signed( -{ 1'b0,x511 } )+$signed( -{ 2'b0,x767 }<<<3'd1 )+$signed(11'd40);
assign y255=temp_y[255][11] ==1'b1 ? 5'd0 :  
        temp_y[255][8] ==1'b1 ? 5'd31 : 
        temp_y[255][2]==1'b1 ? temp_y[255][7:3]+1'b1 : temp_y[255][7:3];
assign temp_y[319] = 
+$signed( -{ 1'b0,x238 } )+$signed( { 2'b0,x494 } <<<3'd1 )+$signed( -{ 1'b0,x750 } )+$signed( -{ 1'b0,x239 } )+$signed( { 2'b0,x495 } <<<3'd1 )+$signed( -{ 2'b0,x751 }<<<3'd1 )+$signed( -{ 1'b0,x254 } )+$signed( { 2'b0,x510 } <<<3'd1 )+$signed( -{ 1'b0,x766 } )+$signed( -{ 2'b0,x255 }<<<3'd1 )+$signed( { 3'b0,x511 }<<<3'd2 )+$signed( -{ 2'b0,x767 }<<<3'd1 )+$signed(11'd32);
assign y319=temp_y[319][11] ==1'b1 ? 5'd0 :  
        temp_y[319][8] ==1'b1 ? 5'd31 : 
        temp_y[319][2]==1'b1 ? temp_y[319][7:3]+1'b1 : temp_y[319][7:3];
assign temp_y[383] = 
+$signed( -{ 1'b0,x238 } )+$signed( -{ 2'b0,x494 }<<<3'd1 )+$signed( -{ 1'b0,x750 } )+$signed( { 1'b0,x239 }  )+$signed( { 2'b0,x495 } <<<3'd1 )+$signed( { 1'b0,x751 }  )+$signed( { 1'b0,x254 }  )+$signed( { 2'b0,x510 } <<<3'd1 )+$signed( { 2'b0,x766 } <<<3'd1 )+$signed( -{ 1'b0,x255 } )+$signed( -{ 2'b0,x511 }<<<3'd1 )+$signed( -{ 1'b0,x767 } )-$signed(11'd68);
assign y383=temp_y[383][11] ==1'b1 ? 5'd0 :  
        temp_y[383][8] ==1'b1 ? 5'd31 : 
        temp_y[383][2]==1'b1 ? temp_y[383][7:3]+1'b1 : temp_y[383][7:3];
assign temp_y[447] = 
+$signed( { 1'b0,x494 }  )+$signed( { 1'b0,x751 }  )+$signed( { 1'b0,x767 }  )-$signed(11'd108);
assign y447=temp_y[447][11] ==1'b1 ? 5'd0 :  
        temp_y[447][8] ==1'b1 ? 5'd31 : 
        temp_y[447][2]==1'b1 ? temp_y[447][7:3]+1'b1 : temp_y[447][7:3];
assign temp_y[511] = 
+$signed( -{ 2'b0,x238 }<<<3'd1 )+$signed( { 2'b0,x750 } <<<3'd1 )+$signed( -{ 2'b0,x239 }<<<3'd1 )+$signed( { 1'b0,x495 }  )+$signed( { 1'b0,x751 }  )+$signed( -{ 2'b0,x254 }<<<3'd1 )+$signed( { 1'b0,x510 }  )+$signed( { 1'b0,x766 }  )+$signed( -{ 1'b0,x255 } )+$signed(11'd64);
assign y511=temp_y[511][11] ==1'b1 ? 5'd0 :  
        temp_y[511][8] ==1'b1 ? 5'd31 : 
        temp_y[511][2]==1'b1 ? temp_y[511][7:3]+1'b1 : temp_y[511][7:3];
assign temp_y[575] = 
+$signed( -{ 2'b0,x238 }<<<3'd1 )+$signed( -{ 1'b0,x494 } )+$signed( -{ 3'b0,x239 }<<<3'd2)+$signed( { 1'b0,x254 }  )+$signed( { 1'b0,x510 }  )+$signed( { 3'b0,x255 }<<<3'd2 )+$signed(11'd16);
assign y575=temp_y[575][11] ==1'b1 ? 5'd0 :  
        temp_y[575][8] ==1'b1 ? 5'd31 : 
        temp_y[575][2]==1'b1 ? temp_y[575][7:3]+1'b1 : temp_y[575][7:3];
assign temp_y[639] = 
+$signed( { 2'b0,x494 } <<<3'd1 )+$signed( { 2'b0,x750 } <<<3'd1 )+$signed( -{ 1'b0,x239 } )+$signed( -{ 2'b0,x495 }<<<3'd1 )+$signed( -{ 2'b0,x751 }<<<3'd1 )+$signed( { 2'b0,x510 } <<<3'd1 )+$signed( { 1'b0,x766 }  )+$signed( -{ 2'b0,x511 }<<<3'd1 )-$signed(11'd8);
assign y639=temp_y[639][11] ==1'b1 ? 5'd0 :  
        temp_y[639][8] ==1'b1 ? 5'd31 : 
        temp_y[639][2]==1'b1 ? temp_y[639][7:3]+1'b1 : temp_y[639][7:3];
endmodule