module top(
input [7:0] x0 ,
input [7:0] x1 ,
input [7:0] x2 ,
input [7:0] x3 ,
input [7:0] x4 ,
input [7:0] x5 ,
input [7:0] x6 ,
input [7:0] x7 ,
input [7:0] x8 ,
input [7:0] x9 ,
input [7:0] x10 ,
input [7:0] x11 ,
input [7:0] x12 ,
input [7:0] x13 ,
input [7:0] x14 ,
input [7:0] x15 ,
input [7:0] x16 ,
input [7:0] x17 ,
input [7:0] x18 ,
input [7:0] x19 ,
input [7:0] x20 ,
input [7:0] x21 ,
input [7:0] x22 ,
input [7:0] x23 ,
input [7:0] x24 ,
input [7:0] x25 ,
input [7:0] x26 ,
input [7:0] x27 ,
input [7:0] x28 ,
input [7:0] x29 ,
input [7:0] x30 ,
input [7:0] x31 ,
input [7:0] x32 ,
input [7:0] x33 ,
input [7:0] x34 ,
input [7:0] x35 ,
input [7:0] x36 ,
input [7:0] x37 ,
input [7:0] x38 ,
input [7:0] x39 ,
input [7:0] x40 ,
input [7:0] x41 ,
input [7:0] x42 ,
input [7:0] x43 ,
input [7:0] x44 ,
input [7:0] x45 ,
input [7:0] x46 ,
input [7:0] x47 ,
input [7:0] x48 ,
input [7:0] x49 ,
input [7:0] x50 ,
input [7:0] x51 ,
input [7:0] x52 ,
input [7:0] x53 ,
input [7:0] x54 ,
input [7:0] x55 ,
input [7:0] x56 ,
input [7:0] x57 ,
input [7:0] x58 ,
input [7:0] x59 ,
input [7:0] x60 ,
input [7:0] x61 ,
input [7:0] x62 ,
input [7:0] x63 ,
input [7:0] x64 ,
input [7:0] x65 ,
input [7:0] x66 ,
input [7:0] x67 ,
input [7:0] x68 ,
input [7:0] x69 ,
input [7:0] x70 ,
input [7:0] x71 ,
input [7:0] x72 ,
input [7:0] x73 ,
input [7:0] x74 ,
input [7:0] x75 ,
input [7:0] x76 ,
input [7:0] x77 ,
input [7:0] x78 ,
input [7:0] x79 ,
input [7:0] x80 ,
input [7:0] x81 ,
input [7:0] x82 ,
input [7:0] x83 ,
input [7:0] x84 ,
input [7:0] x85 ,
input [7:0] x86 ,
input [7:0] x87 ,
input [7:0] x88 ,
input [7:0] x89 ,
input [7:0] x90 ,
input [7:0] x91 ,
input [7:0] x92 ,
input [7:0] x93 ,
input [7:0] x94 ,
input [7:0] x95 ,
input [7:0] x96 ,
input [7:0] x97 ,
input [7:0] x98 ,
input [7:0] x99 ,
input [7:0] x100 ,
input [7:0] x101 ,
input [7:0] x102 ,
input [7:0] x103 ,
input [7:0] x104 ,
input [7:0] x105 ,
input [7:0] x106 ,
input [7:0] x107 ,
input [7:0] x108 ,
input [7:0] x109 ,
input [7:0] x110 ,
input [7:0] x111 ,
input [7:0] x112 ,
input [7:0] x113 ,
input [7:0] x114 ,
input [7:0] x115 ,
input [7:0] x116 ,
input [7:0] x117 ,
input [7:0] x118 ,
input [7:0] x119 ,
input [7:0] x120 ,
input [7:0] x121 ,
input [7:0] x122 ,
input [7:0] x123 ,
input [7:0] x124 ,
input [7:0] x125 ,
input [7:0] x126 ,
input [7:0] x127 ,
input [7:0] x128 ,
input [7:0] x129 ,
input [7:0] x130 ,
input [7:0] x131 ,
input [7:0] x132 ,
input [7:0] x133 ,
input [7:0] x134 ,
input [7:0] x135 ,
input [7:0] x136 ,
input [7:0] x137 ,
input [7:0] x138 ,
input [7:0] x139 ,
input [7:0] x140 ,
input [7:0] x141 ,
input [7:0] x142 ,
input [7:0] x143 ,
input [7:0] x144 ,
input [7:0] x145 ,
input [7:0] x146 ,
input [7:0] x147 ,
input [7:0] x148 ,
input [7:0] x149 ,
input [7:0] x150 ,
input [7:0] x151 ,
input [7:0] x152 ,
input [7:0] x153 ,
input [7:0] x154 ,
input [7:0] x155 ,
input [7:0] x156 ,
input [7:0] x157 ,
input [7:0] x158 ,
input [7:0] x159 ,
input [7:0] x160 ,
input [7:0] x161 ,
input [7:0] x162 ,
input [7:0] x163 ,
input [7:0] x164 ,
input [7:0] x165 ,
input [7:0] x166 ,
input [7:0] x167 ,
input [7:0] x168 ,
input [7:0] x169 ,
input [7:0] x170 ,
input [7:0] x171 ,
input [7:0] x172 ,
input [7:0] x173 ,
input [7:0] x174 ,
input [7:0] x175 ,
input [7:0] x176 ,
input [7:0] x177 ,
input [7:0] x178 ,
input [7:0] x179 ,
input [7:0] x180 ,
input [7:0] x181 ,
input [7:0] x182 ,
input [7:0] x183 ,
input [7:0] x184 ,
input [7:0] x185 ,
input [7:0] x186 ,
input [7:0] x187 ,
input [7:0] x188 ,
input [7:0] x189 ,
input [7:0] x190 ,
input [7:0] x191 ,
input [7:0] x192 ,
input [7:0] x193 ,
input [7:0] x194 ,
input [7:0] x195 ,
input [7:0] x196 ,
input [7:0] x197 ,
input [7:0] x198 ,
input [7:0] x199 ,
input [7:0] x200 ,
input [7:0] x201 ,
input [7:0] x202 ,
input [7:0] x203 ,
input [7:0] x204 ,
input [7:0] x205 ,
input [7:0] x206 ,
input [7:0] x207 ,
input [7:0] x208 ,
input [7:0] x209 ,
input [7:0] x210 ,
input [7:0] x211 ,
input [7:0] x212 ,
input [7:0] x213 ,
input [7:0] x214 ,
input [7:0] x215 ,
input [7:0] x216 ,
input [7:0] x217 ,
input [7:0] x218 ,
input [7:0] x219 ,
input [7:0] x220 ,
input [7:0] x221 ,
input [7:0] x222 ,
input [7:0] x223 ,
input [7:0] x224 ,
input [7:0] x225 ,
input [7:0] x226 ,
input [7:0] x227 ,
input [7:0] x228 ,
input [7:0] x229 ,
input [7:0] x230 ,
input [7:0] x231 ,
input [7:0] x232 ,
input [7:0] x233 ,
input [7:0] x234 ,
input [7:0] x235 ,
input [7:0] x236 ,
input [7:0] x237 ,
input [7:0] x238 ,
input [7:0] x239 ,
input [7:0] x240 ,
input [7:0] x241 ,
input [7:0] x242 ,
input [7:0] x243 ,
input [7:0] x244 ,
input [7:0] x245 ,
input [7:0] x246 ,
input [7:0] x247 ,
input [7:0] x248 ,
input [7:0] x249 ,
input [7:0] x250 ,
input [7:0] x251 ,
input [7:0] x252 ,
input [7:0] x253 ,
input [7:0] x254 ,
input [7:0] x255 ,
input [7:0] x256 ,
input [7:0] x257 ,
input [7:0] x258 ,
input [7:0] x259 ,
input [7:0] x260 ,
input [7:0] x261 ,
input [7:0] x262 ,
input [7:0] x263 ,
input [7:0] x264 ,
input [7:0] x265 ,
input [7:0] x266 ,
input [7:0] x267 ,
input [7:0] x268 ,
input [7:0] x269 ,
input [7:0] x270 ,
input [7:0] x271 ,
input [7:0] x272 ,
input [7:0] x273 ,
input [7:0] x274 ,
input [7:0] x275 ,
input [7:0] x276 ,
input [7:0] x277 ,
input [7:0] x278 ,
input [7:0] x279 ,
input [7:0] x280 ,
input [7:0] x281 ,
input [7:0] x282 ,
input [7:0] x283 ,
input [7:0] x284 ,
input [7:0] x285 ,
input [7:0] x286 ,
input [7:0] x287 ,
input [7:0] x288 ,
input [7:0] x289 ,
input [7:0] x290 ,
input [7:0] x291 ,
input [7:0] x292 ,
input [7:0] x293 ,
input [7:0] x294 ,
input [7:0] x295 ,
input [7:0] x296 ,
input [7:0] x297 ,
input [7:0] x298 ,
input [7:0] x299 ,
input [7:0] x300 ,
input [7:0] x301 ,
input [7:0] x302 ,
input [7:0] x303 ,
input [7:0] x304 ,
input [7:0] x305 ,
input [7:0] x306 ,
input [7:0] x307 ,
input [7:0] x308 ,
input [7:0] x309 ,
input [7:0] x310 ,
input [7:0] x311 ,
input [7:0] x312 ,
input [7:0] x313 ,
input [7:0] x314 ,
input [7:0] x315 ,
input [7:0] x316 ,
input [7:0] x317 ,
input [7:0] x318 ,
input [7:0] x319 ,
input [7:0] x320 ,
input [7:0] x321 ,
input [7:0] x322 ,
input [7:0] x323 ,
input [7:0] x324 ,
input [7:0] x325 ,
input [7:0] x326 ,
input [7:0] x327 ,
input [7:0] x328 ,
input [7:0] x329 ,
input [7:0] x330 ,
input [7:0] x331 ,
input [7:0] x332 ,
input [7:0] x333 ,
input [7:0] x334 ,
input [7:0] x335 ,
input [7:0] x336 ,
input [7:0] x337 ,
input [7:0] x338 ,
input [7:0] x339 ,
input [7:0] x340 ,
input [7:0] x341 ,
input [7:0] x342 ,
input [7:0] x343 ,
input [7:0] x344 ,
input [7:0] x345 ,
input [7:0] x346 ,
input [7:0] x347 ,
input [7:0] x348 ,
input [7:0] x349 ,
input [7:0] x350 ,
input [7:0] x351 ,
input [7:0] x352 ,
input [7:0] x353 ,
input [7:0] x354 ,
input [7:0] x355 ,
input [7:0] x356 ,
input [7:0] x357 ,
input [7:0] x358 ,
input [7:0] x359 ,
input [7:0] x360 ,
input [7:0] x361 ,
input [7:0] x362 ,
input [7:0] x363 ,
input [7:0] x364 ,
input [7:0] x365 ,
input [7:0] x366 ,
input [7:0] x367 ,
input [7:0] x368 ,
input [7:0] x369 ,
input [7:0] x370 ,
input [7:0] x371 ,
input [7:0] x372 ,
input [7:0] x373 ,
input [7:0] x374 ,
input [7:0] x375 ,
input [7:0] x376 ,
input [7:0] x377 ,
input [7:0] x378 ,
input [7:0] x379 ,
input [7:0] x380 ,
input [7:0] x381 ,
input [7:0] x382 ,
input [7:0] x383 ,
input [7:0] x384 ,
input [7:0] x385 ,
input [7:0] x386 ,
input [7:0] x387 ,
input [7:0] x388 ,
input [7:0] x389 ,
input [7:0] x390 ,
input [7:0] x391 ,
input [7:0] x392 ,
input [7:0] x393 ,
input [7:0] x394 ,
input [7:0] x395 ,
input [7:0] x396 ,
input [7:0] x397 ,
input [7:0] x398 ,
input [7:0] x399 ,
input [7:0] x400 ,
input [7:0] x401 ,
input [7:0] x402 ,
input [7:0] x403 ,
input [7:0] x404 ,
input [7:0] x405 ,
input [7:0] x406 ,
input [7:0] x407 ,
input [7:0] x408 ,
input [7:0] x409 ,
input [7:0] x410 ,
input [7:0] x411 ,
input [7:0] x412 ,
input [7:0] x413 ,
input [7:0] x414 ,
input [7:0] x415 ,
input [7:0] x416 ,
input [7:0] x417 ,
input [7:0] x418 ,
input [7:0] x419 ,
input [7:0] x420 ,
input [7:0] x421 ,
input [7:0] x422 ,
input [7:0] x423 ,
input [7:0] x424 ,
input [7:0] x425 ,
input [7:0] x426 ,
input [7:0] x427 ,
input [7:0] x428 ,
input [7:0] x429 ,
input [7:0] x430 ,
input [7:0] x431 ,
input [7:0] x432 ,
input [7:0] x433 ,
input [7:0] x434 ,
input [7:0] x435 ,
input [7:0] x436 ,
input [7:0] x437 ,
input [7:0] x438 ,
input [7:0] x439 ,
input [7:0] x440 ,
input [7:0] x441 ,
input [7:0] x442 ,
input [7:0] x443 ,
input [7:0] x444 ,
input [7:0] x445 ,
input [7:0] x446 ,
input [7:0] x447 ,
input [7:0] x448 ,
input [7:0] x449 ,
input [7:0] x450 ,
input [7:0] x451 ,
input [7:0] x452 ,
input [7:0] x453 ,
input [7:0] x454 ,
input [7:0] x455 ,
input [7:0] x456 ,
input [7:0] x457 ,
input [7:0] x458 ,
input [7:0] x459 ,
input [7:0] x460 ,
input [7:0] x461 ,
input [7:0] x462 ,
input [7:0] x463 ,
input [7:0] x464 ,
input [7:0] x465 ,
input [7:0] x466 ,
input [7:0] x467 ,
input [7:0] x468 ,
input [7:0] x469 ,
input [7:0] x470 ,
input [7:0] x471 ,
input [7:0] x472 ,
input [7:0] x473 ,
input [7:0] x474 ,
input [7:0] x475 ,
input [7:0] x476 ,
input [7:0] x477 ,
input [7:0] x478 ,
input [7:0] x479 ,
input [7:0] x480 ,
input [7:0] x481 ,
input [7:0] x482 ,
input [7:0] x483 ,
input [7:0] x484 ,
input [7:0] x485 ,
input [7:0] x486 ,
input [7:0] x487 ,
input [7:0] x488 ,
input [7:0] x489 ,
input [7:0] x490 ,
input [7:0] x491 ,
input [7:0] x492 ,
input [7:0] x493 ,
input [7:0] x494 ,
input [7:0] x495 ,
input [7:0] x496 ,
input [7:0] x497 ,
input [7:0] x498 ,
input [7:0] x499 ,
input [7:0] x500 ,
input [7:0] x501 ,
input [7:0] x502 ,
input [7:0] x503 ,
input [7:0] x504 ,
input [7:0] x505 ,
input [7:0] x506 ,
input [7:0] x507 ,
input [7:0] x508 ,
input [7:0] x509 ,
input [7:0] x510 ,
input [7:0] x511 ,
input [7:0] x512 ,
input [7:0] x513 ,
input [7:0] x514 ,
input [7:0] x515 ,
input [7:0] x516 ,
input [7:0] x517 ,
input [7:0] x518 ,
input [7:0] x519 ,
input [7:0] x520 ,
input [7:0] x521 ,
input [7:0] x522 ,
input [7:0] x523 ,
input [7:0] x524 ,
input [7:0] x525 ,
input [7:0] x526 ,
input [7:0] x527 ,
input [7:0] x528 ,
input [7:0] x529 ,
input [7:0] x530 ,
input [7:0] x531 ,
input [7:0] x532 ,
input [7:0] x533 ,
input [7:0] x534 ,
input [7:0] x535 ,
input [7:0] x536 ,
input [7:0] x537 ,
input [7:0] x538 ,
input [7:0] x539 ,
input [7:0] x540 ,
input [7:0] x541 ,
input [7:0] x542 ,
input [7:0] x543 ,
input [7:0] x544 ,
input [7:0] x545 ,
input [7:0] x546 ,
input [7:0] x547 ,
input [7:0] x548 ,
input [7:0] x549 ,
input [7:0] x550 ,
input [7:0] x551 ,
input [7:0] x552 ,
input [7:0] x553 ,
input [7:0] x554 ,
input [7:0] x555 ,
input [7:0] x556 ,
input [7:0] x557 ,
input [7:0] x558 ,
input [7:0] x559 ,
input [7:0] x560 ,
input [7:0] x561 ,
input [7:0] x562 ,
input [7:0] x563 ,
input [7:0] x564 ,
input [7:0] x565 ,
input [7:0] x566 ,
input [7:0] x567 ,
input [7:0] x568 ,
input [7:0] x569 ,
input [7:0] x570 ,
input [7:0] x571 ,
input [7:0] x572 ,
input [7:0] x573 ,
input [7:0] x574 ,
input [7:0] x575 ,
input [7:0] x576 ,
input [7:0] x577 ,
input [7:0] x578 ,
input [7:0] x579 ,
input [7:0] x580 ,
input [7:0] x581 ,
input [7:0] x582 ,
input [7:0] x583 ,
input [7:0] x584 ,
input [7:0] x585 ,
input [7:0] x586 ,
input [7:0] x587 ,
input [7:0] x588 ,
input [7:0] x589 ,
input [7:0] x590 ,
input [7:0] x591 ,
input [7:0] x592 ,
input [7:0] x593 ,
input [7:0] x594 ,
input [7:0] x595 ,
input [7:0] x596 ,
input [7:0] x597 ,
input [7:0] x598 ,
input [7:0] x599 ,
input [7:0] x600 ,
input [7:0] x601 ,
input [7:0] x602 ,
input [7:0] x603 ,
input [7:0] x604 ,
input [7:0] x605 ,
input [7:0] x606 ,
input [7:0] x607 ,
input [7:0] x608 ,
input [7:0] x609 ,
input [7:0] x610 ,
input [7:0] x611 ,
input [7:0] x612 ,
input [7:0] x613 ,
input [7:0] x614 ,
input [7:0] x615 ,
input [7:0] x616 ,
input [7:0] x617 ,
input [7:0] x618 ,
input [7:0] x619 ,
input [7:0] x620 ,
input [7:0] x621 ,
input [7:0] x622 ,
input [7:0] x623 ,
input [7:0] x624 ,
input [7:0] x625 ,
input [7:0] x626 ,
input [7:0] x627 ,
input [7:0] x628 ,
input [7:0] x629 ,
input [7:0] x630 ,
input [7:0] x631 ,
input [7:0] x632 ,
input [7:0] x633 ,
input [7:0] x634 ,
input [7:0] x635 ,
input [7:0] x636 ,
input [7:0] x637 ,
input [7:0] x638 ,
input [7:0] x639 ,
input [7:0] x640 ,
input [7:0] x641 ,
input [7:0] x642 ,
input [7:0] x643 ,
input [7:0] x644 ,
input [7:0] x645 ,
input [7:0] x646 ,
input [7:0] x647 ,
input [7:0] x648 ,
input [7:0] x649 ,
input [7:0] x650 ,
input [7:0] x651 ,
input [7:0] x652 ,
input [7:0] x653 ,
input [7:0] x654 ,
input [7:0] x655 ,
input [7:0] x656 ,
input [7:0] x657 ,
input [7:0] x658 ,
input [7:0] x659 ,
input [7:0] x660 ,
input [7:0] x661 ,
input [7:0] x662 ,
input [7:0] x663 ,
input [7:0] x664 ,
input [7:0] x665 ,
input [7:0] x666 ,
input [7:0] x667 ,
input [7:0] x668 ,
input [7:0] x669 ,
input [7:0] x670 ,
input [7:0] x671 ,
input [7:0] x672 ,
input [7:0] x673 ,
input [7:0] x674 ,
input [7:0] x675 ,
input [7:0] x676 ,
input [7:0] x677 ,
input [7:0] x678 ,
input [7:0] x679 ,
input [7:0] x680 ,
input [7:0] x681 ,
input [7:0] x682 ,
input [7:0] x683 ,
input [7:0] x684 ,
input [7:0] x685 ,
input [7:0] x686 ,
input [7:0] x687 ,
input [7:0] x688 ,
input [7:0] x689 ,
input [7:0] x690 ,
input [7:0] x691 ,
input [7:0] x692 ,
input [7:0] x693 ,
input [7:0] x694 ,
input [7:0] x695 ,
input [7:0] x696 ,
input [7:0] x697 ,
input [7:0] x698 ,
input [7:0] x699 ,
input [7:0] x700 ,
input [7:0] x701 ,
input [7:0] x702 ,
input [7:0] x703 ,
input [7:0] x704 ,
input [7:0] x705 ,
input [7:0] x706 ,
input [7:0] x707 ,
input [7:0] x708 ,
input [7:0] x709 ,
input [7:0] x710 ,
input [7:0] x711 ,
input [7:0] x712 ,
input [7:0] x713 ,
input [7:0] x714 ,
input [7:0] x715 ,
input [7:0] x716 ,
input [7:0] x717 ,
input [7:0] x718 ,
input [7:0] x719 ,
input [7:0] x720 ,
input [7:0] x721 ,
input [7:0] x722 ,
input [7:0] x723 ,
input [7:0] x724 ,
input [7:0] x725 ,
input [7:0] x726 ,
input [7:0] x727 ,
input [7:0] x728 ,
input [7:0] x729 ,
input [7:0] x730 ,
input [7:0] x731 ,
input [7:0] x732 ,
input [7:0] x733 ,
input [7:0] x734 ,
input [7:0] x735 ,
input [7:0] x736 ,
input [7:0] x737 ,
input [7:0] x738 ,
input [7:0] x739 ,
input [7:0] x740 ,
input [7:0] x741 ,
input [7:0] x742 ,
input [7:0] x743 ,
input [7:0] x744 ,
input [7:0] x745 ,
input [7:0] x746 ,
input [7:0] x747 ,
input [7:0] x748 ,
input [7:0] x749 ,
input [7:0] x750 ,
input [7:0] x751 ,
input [7:0] x752 ,
input [7:0] x753 ,
input [7:0] x754 ,
input [7:0] x755 ,
input [7:0] x756 ,
input [7:0] x757 ,
input [7:0] x758 ,
input [7:0] x759 ,
input [7:0] x760 ,
input [7:0] x761 ,
input [7:0] x762 ,
input [7:0] x763 ,
input [7:0] x764 ,
input [7:0] x765 ,
input [7:0] x766 ,
input [7:0] x767 ,
input [7:0] x768 ,
input [7:0] x769 ,
input [7:0] x770 ,
input [7:0] x771 ,
input [7:0] x772 ,
input [7:0] x773 ,
input [7:0] x774 ,
input [7:0] x775 ,
input [7:0] x776 ,
input [7:0] x777 ,
input [7:0] x778 ,
input [7:0] x779 ,
input [7:0] x780 ,
input [7:0] x781 ,
input [7:0] x782 ,
input [7:0] x783 ,
input [7:0] x784 ,
input [7:0] x785 ,
input [7:0] x786 ,
input [7:0] x787 ,
input [7:0] x788 ,
input [7:0] x789 ,
input [7:0] x790 ,
input [7:0] x791 ,
input [7:0] x792 ,
input [7:0] x793 ,
input [7:0] x794 ,
input [7:0] x795 ,
input [7:0] x796 ,
input [7:0] x797 ,
input [7:0] x798 ,
input [7:0] x799 ,
input [7:0] x800 ,
input [7:0] x801 ,
input [7:0] x802 ,
input [7:0] x803 ,
input [7:0] x804 ,
input [7:0] x805 ,
input [7:0] x806 ,
input [7:0] x807 ,
input [7:0] x808 ,
input [7:0] x809 ,
input [7:0] x810 ,
input [7:0] x811 ,
input [7:0] x812 ,
input [7:0] x813 ,
input [7:0] x814 ,
input [7:0] x815 ,
input [7:0] x816 ,
input [7:0] x817 ,
input [7:0] x818 ,
input [7:0] x819 ,
input [7:0] x820 ,
input [7:0] x821 ,
input [7:0] x822 ,
input [7:0] x823 ,
input [7:0] x824 ,
input [7:0] x825 ,
input [7:0] x826 ,
input [7:0] x827 ,
input [7:0] x828 ,
input [7:0] x829 ,
input [7:0] x830 ,
input [7:0] x831 ,
input [7:0] x832 ,
input [7:0] x833 ,
input [7:0] x834 ,
input [7:0] x835 ,
input [7:0] x836 ,
input [7:0] x837 ,
input [7:0] x838 ,
input [7:0] x839 ,
input [7:0] x840 ,
input [7:0] x841 ,
input [7:0] x842 ,
input [7:0] x843 ,
input [7:0] x844 ,
input [7:0] x845 ,
input [7:0] x846 ,
input [7:0] x847 ,
input [7:0] x848 ,
input [7:0] x849 ,
input [7:0] x850 ,
input [7:0] x851 ,
input [7:0] x852 ,
input [7:0] x853 ,
input [7:0] x854 ,
input [7:0] x855 ,
input [7:0] x856 ,
input [7:0] x857 ,
input [7:0] x858 ,
input [7:0] x859 ,
input [7:0] x860 ,
input [7:0] x861 ,
input [7:0] x862 ,
input [7:0] x863 ,
input [7:0] x864 ,
input [7:0] x865 ,
input [7:0] x866 ,
input [7:0] x867 ,
input [7:0] x868 ,
input [7:0] x869 ,
input [7:0] x870 ,
input [7:0] x871 ,
input [7:0] x872 ,
input [7:0] x873 ,
input [7:0] x874 ,
input [7:0] x875 ,
input [7:0] x876 ,
input [7:0] x877 ,
input [7:0] x878 ,
input [7:0] x879 ,
input [7:0] x880 ,
input [7:0] x881 ,
input [7:0] x882 ,
input [7:0] x883 ,
input [7:0] x884 ,
input [7:0] x885 ,
input [7:0] x886 ,
input [7:0] x887 ,
input [7:0] x888 ,
input [7:0] x889 ,
input [7:0] x890 ,
input [7:0] x891 ,
input [7:0] x892 ,
input [7:0] x893 ,
input [7:0] x894 ,
input [7:0] x895 ,
input [7:0] x896 ,
input [7:0] x897 ,
input [7:0] x898 ,
input [7:0] x899 ,
input [7:0] x900 ,
input [7:0] x901 ,
input [7:0] x902 ,
input [7:0] x903 ,
input [7:0] x904 ,
input [7:0] x905 ,
input [7:0] x906 ,
input [7:0] x907 ,
input [7:0] x908 ,
input [7:0] x909 ,
input [7:0] x910 ,
input [7:0] x911 ,
input [7:0] x912 ,
input [7:0] x913 ,
input [7:0] x914 ,
input [7:0] x915 ,
input [7:0] x916 ,
input [7:0] x917 ,
input [7:0] x918 ,
input [7:0] x919 ,
input [7:0] x920 ,
input [7:0] x921 ,
input [7:0] x922 ,
input [7:0] x923 ,
input [7:0] x924 ,
input [7:0] x925 ,
input [7:0] x926 ,
input [7:0] x927 ,
input [7:0] x928 ,
input [7:0] x929 ,
input [7:0] x930 ,
input [7:0] x931 ,
input [7:0] x932 ,
input [7:0] x933 ,
input [7:0] x934 ,
input [7:0] x935 ,
input [7:0] x936 ,
input [7:0] x937 ,
input [7:0] x938 ,
input [7:0] x939 ,
input [7:0] x940 ,
input [7:0] x941 ,
input [7:0] x942 ,
input [7:0] x943 ,
input [7:0] x944 ,
input [7:0] x945 ,
input [7:0] x946 ,
input [7:0] x947 ,
input [7:0] x948 ,
input [7:0] x949 ,
input [7:0] x950 ,
input [7:0] x951 ,
input [7:0] x952 ,
input [7:0] x953 ,
input [7:0] x954 ,
input [7:0] x955 ,
input [7:0] x956 ,
input [7:0] x957 ,
input [7:0] x958 ,
input [7:0] x959 ,
input [7:0] x960 ,
input [7:0] x961 ,
input [7:0] x962 ,
input [7:0] x963 ,
input [7:0] x964 ,
input [7:0] x965 ,
input [7:0] x966 ,
input [7:0] x967 ,
input [7:0] x968 ,
input [7:0] x969 ,
input [7:0] x970 ,
input [7:0] x971 ,
input [7:0] x972 ,
input [7:0] x973 ,
input [7:0] x974 ,
input [7:0] x975 ,
input [7:0] x976 ,
input [7:0] x977 ,
input [7:0] x978 ,
input [7:0] x979 ,
input [7:0] x980 ,
input [7:0] x981 ,
input [7:0] x982 ,
input [7:0] x983 ,
input [7:0] x984 ,
input [7:0] x985 ,
input [7:0] x986 ,
input [7:0] x987 ,
input [7:0] x988 ,
input [7:0] x989 ,
input [7:0] x990 ,
input [7:0] x991 ,
input [7:0] x992 ,
input [7:0] x993 ,
input [7:0] x994 ,
input [7:0] x995 ,
input [7:0] x996 ,
input [7:0] x997 ,
input [7:0] x998 ,
input [7:0] x999 ,
input [7:0] x1000 ,
input [7:0] x1001 ,
input [7:0] x1002 ,
input [7:0] x1003 ,
input [7:0] x1004 ,
input [7:0] x1005 ,
input [7:0] x1006 ,
input [7:0] x1007 ,
input [7:0] x1008 ,
input [7:0] x1009 ,
input [7:0] x1010 ,
input [7:0] x1011 ,
input [7:0] x1012 ,
input [7:0] x1013 ,
input [7:0] x1014 ,
input [7:0] x1015 ,
input [7:0] x1016 ,
input [7:0] x1017 ,
input [7:0] x1018 ,
input [7:0] x1019 ,
input [7:0] x1020 ,
input [7:0] x1021 ,
input [7:0] x1022 ,
input [7:0] x1023 ,
input [7:0] x1024 ,
input [7:0] x1025 ,
input [7:0] x1026 ,
input [7:0] x1027 ,
input [7:0] x1028 ,
input [7:0] x1029 ,
input [7:0] x1030 ,
input [7:0] x1031 ,
input [7:0] x1032 ,
input [7:0] x1033 ,
input [7:0] x1034 ,
input [7:0] x1035 ,
input [7:0] x1036 ,
input [7:0] x1037 ,
input [7:0] x1038 ,
input [7:0] x1039 ,
input [7:0] x1040 ,
input [7:0] x1041 ,
input [7:0] x1042 ,
input [7:0] x1043 ,
input [7:0] x1044 ,
input [7:0] x1045 ,
input [7:0] x1046 ,
input [7:0] x1047 ,
input [7:0] x1048 ,
input [7:0] x1049 ,
input [7:0] x1050 ,
input [7:0] x1051 ,
input [7:0] x1052 ,
input [7:0] x1053 ,
input [7:0] x1054 ,
input [7:0] x1055 ,
input [7:0] x1056 ,
input [7:0] x1057 ,
input [7:0] x1058 ,
input [7:0] x1059 ,
input [7:0] x1060 ,
input [7:0] x1061 ,
input [7:0] x1062 ,
input [7:0] x1063 ,
input [7:0] x1064 ,
input [7:0] x1065 ,
input [7:0] x1066 ,
input [7:0] x1067 ,
input [7:0] x1068 ,
input [7:0] x1069 ,
input [7:0] x1070 ,
input [7:0] x1071 ,
input [7:0] x1072 ,
input [7:0] x1073 ,
input [7:0] x1074 ,
input [7:0] x1075 ,
input [7:0] x1076 ,
input [7:0] x1077 ,
input [7:0] x1078 ,
input [7:0] x1079 ,
input [7:0] x1080 ,
input [7:0] x1081 ,
input [7:0] x1082 ,
input [7:0] x1083 ,
input [7:0] x1084 ,
input [7:0] x1085 ,
input [7:0] x1086 ,
input [7:0] x1087 ,
input [7:0] x1088 ,
input [7:0] x1089 ,
input [7:0] x1090 ,
input [7:0] x1091 ,
input [7:0] x1092 ,
input [7:0] x1093 ,
input [7:0] x1094 ,
input [7:0] x1095 ,
input [7:0] x1096 ,
input [7:0] x1097 ,
input [7:0] x1098 ,
input [7:0] x1099 ,
input [7:0] x1100 ,
input [7:0] x1101 ,
input [7:0] x1102 ,
input [7:0] x1103 ,
input [7:0] x1104 ,
input [7:0] x1105 ,
input [7:0] x1106 ,
input [7:0] x1107 ,
input [7:0] x1108 ,
input [7:0] x1109 ,
input [7:0] x1110 ,
input [7:0] x1111 ,
input [7:0] x1112 ,
input [7:0] x1113 ,
input [7:0] x1114 ,
input [7:0] x1115 ,
input [7:0] x1116 ,
input [7:0] x1117 ,
input [7:0] x1118 ,
input [7:0] x1119 ,
input [7:0] x1120 ,
input [7:0] x1121 ,
input [7:0] x1122 ,
input [7:0] x1123 ,
input [7:0] x1124 ,
input [7:0] x1125 ,
input [7:0] x1126 ,
input [7:0] x1127 ,
input [7:0] x1128 ,
input [7:0] x1129 ,
input [7:0] x1130 ,
input [7:0] x1131 ,
input [7:0] x1132 ,
input [7:0] x1133 ,
input [7:0] x1134 ,
input [7:0] x1135 ,
input [7:0] x1136 ,
input [7:0] x1137 ,
input [7:0] x1138 ,
input [7:0] x1139 ,
input [7:0] x1140 ,
input [7:0] x1141 ,
input [7:0] x1142 ,
input [7:0] x1143 ,
input [7:0] x1144 ,
input [7:0] x1145 ,
input [7:0] x1146 ,
input [7:0] x1147 ,
input [7:0] x1148 ,
input [7:0] x1149 ,
input [7:0] x1150 ,
input [7:0] x1151 ,
input [7:0] x1152 ,
input [7:0] x1153 ,
input [7:0] x1154 ,
input [7:0] x1155 ,
input [7:0] x1156 ,
input [7:0] x1157 ,
input [7:0] x1158 ,
input [7:0] x1159 ,
input [7:0] x1160 ,
input [7:0] x1161 ,
input [7:0] x1162 ,
input [7:0] x1163 ,
input [7:0] x1164 ,
input [7:0] x1165 ,
input [7:0] x1166 ,
input [7:0] x1167 ,
input [7:0] x1168 ,
input [7:0] x1169 ,
input [7:0] x1170 ,
input [7:0] x1171 ,
input [7:0] x1172 ,
input [7:0] x1173 ,
input [7:0] x1174 ,
input [7:0] x1175 ,
input [7:0] x1176 ,
input [7:0] x1177 ,
input [7:0] x1178 ,
input [7:0] x1179 ,
input [7:0] x1180 ,
input [7:0] x1181 ,
input [7:0] x1182 ,
input [7:0] x1183 ,
input [7:0] x1184 ,
input [7:0] x1185 ,
input [7:0] x1186 ,
input [7:0] x1187 ,
input [7:0] x1188 ,
input [7:0] x1189 ,
input [7:0] x1190 ,
input [7:0] x1191 ,
input [7:0] x1192 ,
input [7:0] x1193 ,
input [7:0] x1194 ,
input [7:0] x1195 ,
input [7:0] x1196 ,
input [7:0] x1197 ,
input [7:0] x1198 ,
input [7:0] x1199 ,
input [7:0] x1200 ,
input [7:0] x1201 ,
input [7:0] x1202 ,
input [7:0] x1203 ,
input [7:0] x1204 ,
input [7:0] x1205 ,
input [7:0] x1206 ,
input [7:0] x1207 ,
input [7:0] x1208 ,
input [7:0] x1209 ,
input [7:0] x1210 ,
input [7:0] x1211 ,
input [7:0] x1212 ,
input [7:0] x1213 ,
input [7:0] x1214 ,
input [7:0] x1215 ,
input [7:0] x1216 ,
input [7:0] x1217 ,
input [7:0] x1218 ,
input [7:0] x1219 ,
input [7:0] x1220 ,
input [7:0] x1221 ,
input [7:0] x1222 ,
input [7:0] x1223 ,
input [7:0] x1224 ,
input [7:0] x1225 ,
input [7:0] x1226 ,
input [7:0] x1227 ,
input [7:0] x1228 ,
input [7:0] x1229 ,
input [7:0] x1230 ,
input [7:0] x1231 ,
input [7:0] x1232 ,
input [7:0] x1233 ,
input [7:0] x1234 ,
input [7:0] x1235 ,
input [7:0] x1236 ,
input [7:0] x1237 ,
input [7:0] x1238 ,
input [7:0] x1239 ,
input [7:0] x1240 ,
input [7:0] x1241 ,
input [7:0] x1242 ,
input [7:0] x1243 ,
input [7:0] x1244 ,
input [7:0] x1245 ,
input [7:0] x1246 ,
input [7:0] x1247 ,
input [7:0] x1248 ,
input [7:0] x1249 ,
input [7:0] x1250 ,
input [7:0] x1251 ,
input [7:0] x1252 ,
input [7:0] x1253 ,
input [7:0] x1254 ,
input [7:0] x1255 ,
input [7:0] x1256 ,
input [7:0] x1257 ,
input [7:0] x1258 ,
input [7:0] x1259 ,
input [7:0] x1260 ,
input [7:0] x1261 ,
input [7:0] x1262 ,
input [7:0] x1263 ,
input [7:0] x1264 ,
input [7:0] x1265 ,
input [7:0] x1266 ,
input [7:0] x1267 ,
input [7:0] x1268 ,
input [7:0] x1269 ,
input [7:0] x1270 ,
input [7:0] x1271 ,
input [7:0] x1272 ,
input [7:0] x1273 ,
input [7:0] x1274 ,
input [7:0] x1275 ,
input [7:0] x1276 ,
input [7:0] x1277 ,
input [7:0] x1278 ,
input [7:0] x1279 ,
input [7:0] x1280 ,
input [7:0] x1281 ,
input [7:0] x1282 ,
input [7:0] x1283 ,
input [7:0] x1284 ,
input [7:0] x1285 ,
input [7:0] x1286 ,
input [7:0] x1287 ,
input [7:0] x1288 ,
input [7:0] x1289 ,
input [7:0] x1290 ,
input [7:0] x1291 ,
input [7:0] x1292 ,
input [7:0] x1293 ,
input [7:0] x1294 ,
input [7:0] x1295 ,
input [7:0] x1296 ,
input [7:0] x1297 ,
input [7:0] x1298 ,
input [7:0] x1299 ,
input [7:0] x1300 ,
input [7:0] x1301 ,
input [7:0] x1302 ,
input [7:0] x1303 ,
input [7:0] x1304 ,
input [7:0] x1305 ,
input [7:0] x1306 ,
input [7:0] x1307 ,
input [7:0] x1308 ,
input [7:0] x1309 ,
input [7:0] x1310 ,
input [7:0] x1311 ,
input [7:0] x1312 ,
input [7:0] x1313 ,
input [7:0] x1314 ,
input [7:0] x1315 ,
input [7:0] x1316 ,
input [7:0] x1317 ,
input [7:0] x1318 ,
input [7:0] x1319 ,
input [7:0] x1320 ,
input [7:0] x1321 ,
input [7:0] x1322 ,
input [7:0] x1323 ,
input [7:0] x1324 ,
input [7:0] x1325 ,
input [7:0] x1326 ,
input [7:0] x1327 ,
input [7:0] x1328 ,
input [7:0] x1329 ,
input [7:0] x1330 ,
input [7:0] x1331 ,
input [7:0] x1332 ,
input [7:0] x1333 ,
input [7:0] x1334 ,
input [7:0] x1335 ,
input [7:0] x1336 ,
input [7:0] x1337 ,
input [7:0] x1338 ,
input [7:0] x1339 ,
input [7:0] x1340 ,
input [7:0] x1341 ,
input [7:0] x1342 ,
input [7:0] x1343 ,
input [7:0] x1344 ,
input [7:0] x1345 ,
input [7:0] x1346 ,
input [7:0] x1347 ,
input [7:0] x1348 ,
input [7:0] x1349 ,
input [7:0] x1350 ,
input [7:0] x1351 ,
input [7:0] x1352 ,
input [7:0] x1353 ,
input [7:0] x1354 ,
input [7:0] x1355 ,
input [7:0] x1356 ,
input [7:0] x1357 ,
input [7:0] x1358 ,
input [7:0] x1359 ,
input [7:0] x1360 ,
input [7:0] x1361 ,
input [7:0] x1362 ,
input [7:0] x1363 ,
input [7:0] x1364 ,
input [7:0] x1365 ,
input [7:0] x1366 ,
input [7:0] x1367 ,
input [7:0] x1368 ,
input [7:0] x1369 ,
input [7:0] x1370 ,
input [7:0] x1371 ,
input [7:0] x1372 ,
input [7:0] x1373 ,
input [7:0] x1374 ,
input [7:0] x1375 ,
input [7:0] x1376 ,
input [7:0] x1377 ,
input [7:0] x1378 ,
input [7:0] x1379 ,
input [7:0] x1380 ,
input [7:0] x1381 ,
input [7:0] x1382 ,
input [7:0] x1383 ,
input [7:0] x1384 ,
input [7:0] x1385 ,
input [7:0] x1386 ,
input [7:0] x1387 ,
input [7:0] x1388 ,
input [7:0] x1389 ,
input [7:0] x1390 ,
input [7:0] x1391 ,
input [7:0] x1392 ,
input [7:0] x1393 ,
input [7:0] x1394 ,
input [7:0] x1395 ,
input [7:0] x1396 ,
input [7:0] x1397 ,
input [7:0] x1398 ,
input [7:0] x1399 ,
input [7:0] x1400 ,
input [7:0] x1401 ,
input [7:0] x1402 ,
input [7:0] x1403 ,
input [7:0] x1404 ,
input [7:0] x1405 ,
input [7:0] x1406 ,
input [7:0] x1407 ,
input [7:0] x1408 ,
input [7:0] x1409 ,
input [7:0] x1410 ,
input [7:0] x1411 ,
input [7:0] x1412 ,
input [7:0] x1413 ,
input [7:0] x1414 ,
input [7:0] x1415 ,
input [7:0] x1416 ,
input [7:0] x1417 ,
input [7:0] x1418 ,
input [7:0] x1419 ,
input [7:0] x1420 ,
input [7:0] x1421 ,
input [7:0] x1422 ,
input [7:0] x1423 ,
input [7:0] x1424 ,
input [7:0] x1425 ,
input [7:0] x1426 ,
input [7:0] x1427 ,
input [7:0] x1428 ,
input [7:0] x1429 ,
input [7:0] x1430 ,
input [7:0] x1431 ,
input [7:0] x1432 ,
input [7:0] x1433 ,
input [7:0] x1434 ,
input [7:0] x1435 ,
input [7:0] x1436 ,
input [7:0] x1437 ,
input [7:0] x1438 ,
input [7:0] x1439 ,
input [7:0] x1440 ,
input [7:0] x1441 ,
input [7:0] x1442 ,
input [7:0] x1443 ,
input [7:0] x1444 ,
input [7:0] x1445 ,
input [7:0] x1446 ,
input [7:0] x1447 ,
input [7:0] x1448 ,
input [7:0] x1449 ,
input [7:0] x1450 ,
input [7:0] x1451 ,
input [7:0] x1452 ,
input [7:0] x1453 ,
input [7:0] x1454 ,
input [7:0] x1455 ,
input [7:0] x1456 ,
input [7:0] x1457 ,
input [7:0] x1458 ,
input [7:0] x1459 ,
input [7:0] x1460 ,
input [7:0] x1461 ,
input [7:0] x1462 ,
input [7:0] x1463 ,
input [7:0] x1464 ,
input [7:0] x1465 ,
input [7:0] x1466 ,
input [7:0] x1467 ,
input [7:0] x1468 ,
input [7:0] x1469 ,
input [7:0] x1470 ,
input [7:0] x1471 ,
input [7:0] x1472 ,
input [7:0] x1473 ,
input [7:0] x1474 ,
input [7:0] x1475 ,
input [7:0] x1476 ,
input [7:0] x1477 ,
input [7:0] x1478 ,
input [7:0] x1479 ,
input [7:0] x1480 ,
input [7:0] x1481 ,
input [7:0] x1482 ,
input [7:0] x1483 ,
input [7:0] x1484 ,
input [7:0] x1485 ,
input [7:0] x1486 ,
input [7:0] x1487 ,
input [7:0] x1488 ,
input [7:0] x1489 ,
input [7:0] x1490 ,
input [7:0] x1491 ,
input [7:0] x1492 ,
input [7:0] x1493 ,
input [7:0] x1494 ,
input [7:0] x1495 ,
input [7:0] x1496 ,
input [7:0] x1497 ,
input [7:0] x1498 ,
input [7:0] x1499 ,
input [7:0] x1500 ,
input [7:0] x1501 ,
input [7:0] x1502 ,
input [7:0] x1503 ,
input [7:0] x1504 ,
input [7:0] x1505 ,
input [7:0] x1506 ,
input [7:0] x1507 ,
input [7:0] x1508 ,
input [7:0] x1509 ,
input [7:0] x1510 ,
input [7:0] x1511 ,
input [7:0] x1512 ,
input [7:0] x1513 ,
input [7:0] x1514 ,
input [7:0] x1515 ,
input [7:0] x1516 ,
input [7:0] x1517 ,
input [7:0] x1518 ,
input [7:0] x1519 ,
input [7:0] x1520 ,
input [7:0] x1521 ,
input [7:0] x1522 ,
input [7:0] x1523 ,
input [7:0] x1524 ,
input [7:0] x1525 ,
input [7:0] x1526 ,
input [7:0] x1527 ,
input [7:0] x1528 ,
input [7:0] x1529 ,
input [7:0] x1530 ,
input [7:0] x1531 ,
input [7:0] x1532 ,
input [7:0] x1533 ,
input [7:0] x1534 ,
input [7:0] x1535 ,
input [7:0] x1536 ,
input [7:0] x1537 ,
input [7:0] x1538 ,
input [7:0] x1539 ,
input [7:0] x1540 ,
input [7:0] x1541 ,
input [7:0] x1542 ,
input [7:0] x1543 ,
input [7:0] x1544 ,
input [7:0] x1545 ,
input [7:0] x1546 ,
input [7:0] x1547 ,
input [7:0] x1548 ,
input [7:0] x1549 ,
input [7:0] x1550 ,
input [7:0] x1551 ,
input [7:0] x1552 ,
input [7:0] x1553 ,
input [7:0] x1554 ,
input [7:0] x1555 ,
input [7:0] x1556 ,
input [7:0] x1557 ,
input [7:0] x1558 ,
input [7:0] x1559 ,
input [7:0] x1560 ,
input [7:0] x1561 ,
input [7:0] x1562 ,
input [7:0] x1563 ,
input [7:0] x1564 ,
input [7:0] x1565 ,
input [7:0] x1566 ,
input [7:0] x1567 ,
input [7:0] x1568 ,
input [7:0] x1569 ,
input [7:0] x1570 ,
input [7:0] x1571 ,
input [7:0] x1572 ,
input [7:0] x1573 ,
input [7:0] x1574 ,
input [7:0] x1575 ,
input [7:0] x1576 ,
input [7:0] x1577 ,
input [7:0] x1578 ,
input [7:0] x1579 ,
input [7:0] x1580 ,
input [7:0] x1581 ,
input [7:0] x1582 ,
input [7:0] x1583 ,
input [7:0] x1584 ,
input [7:0] x1585 ,
input [7:0] x1586 ,
input [7:0] x1587 ,
input [7:0] x1588 ,
input [7:0] x1589 ,
input [7:0] x1590 ,
input [7:0] x1591 ,
input [7:0] x1592 ,
input [7:0] x1593 ,
input [7:0] x1594 ,
input [7:0] x1595 ,
input [7:0] x1596 ,
input [7:0] x1597 ,
input [7:0] x1598 ,
input [7:0] x1599 ,
input [7:0] x1600 ,
input [7:0] x1601 ,
input [7:0] x1602 ,
input [7:0] x1603 ,
input [7:0] x1604 ,
input [7:0] x1605 ,
input [7:0] x1606 ,
input [7:0] x1607 ,
input [7:0] x1608 ,
input [7:0] x1609 ,
input [7:0] x1610 ,
input [7:0] x1611 ,
input [7:0] x1612 ,
input [7:0] x1613 ,
input [7:0] x1614 ,
input [7:0] x1615 ,
input [7:0] x1616 ,
input [7:0] x1617 ,
input [7:0] x1618 ,
input [7:0] x1619 ,
input [7:0] x1620 ,
input [7:0] x1621 ,
input [7:0] x1622 ,
input [7:0] x1623 ,
input [7:0] x1624 ,
input [7:0] x1625 ,
input [7:0] x1626 ,
input [7:0] x1627 ,
input [7:0] x1628 ,
input [7:0] x1629 ,
input [7:0] x1630 ,
input [7:0] x1631 ,
input [7:0] x1632 ,
input [7:0] x1633 ,
input [7:0] x1634 ,
input [7:0] x1635 ,
input [7:0] x1636 ,
input [7:0] x1637 ,
input [7:0] x1638 ,
input [7:0] x1639 ,
input [7:0] x1640 ,
input [7:0] x1641 ,
input [7:0] x1642 ,
input [7:0] x1643 ,
input [7:0] x1644 ,
input [7:0] x1645 ,
input [7:0] x1646 ,
input [7:0] x1647 ,
input [7:0] x1648 ,
input [7:0] x1649 ,
input [7:0] x1650 ,
input [7:0] x1651 ,
input [7:0] x1652 ,
input [7:0] x1653 ,
input [7:0] x1654 ,
input [7:0] x1655 ,
input [7:0] x1656 ,
input [7:0] x1657 ,
input [7:0] x1658 ,
input [7:0] x1659 ,
input [7:0] x1660 ,
input [7:0] x1661 ,
input [7:0] x1662 ,
input [7:0] x1663 ,
input [7:0] x1664 ,
input [7:0] x1665 ,
input [7:0] x1666 ,
input [7:0] x1667 ,
input [7:0] x1668 ,
input [7:0] x1669 ,
input [7:0] x1670 ,
input [7:0] x1671 ,
input [7:0] x1672 ,
input [7:0] x1673 ,
input [7:0] x1674 ,
input [7:0] x1675 ,
input [7:0] x1676 ,
input [7:0] x1677 ,
input [7:0] x1678 ,
input [7:0] x1679 ,
input [7:0] x1680 ,
input [7:0] x1681 ,
input [7:0] x1682 ,
input [7:0] x1683 ,
input [7:0] x1684 ,
input [7:0] x1685 ,
input [7:0] x1686 ,
input [7:0] x1687 ,
input [7:0] x1688 ,
input [7:0] x1689 ,
input [7:0] x1690 ,
input [7:0] x1691 ,
input [7:0] x1692 ,
input [7:0] x1693 ,
input [7:0] x1694 ,
input [7:0] x1695 ,
input [7:0] x1696 ,
input [7:0] x1697 ,
input [7:0] x1698 ,
input [7:0] x1699 ,
input [7:0] x1700 ,
input [7:0] x1701 ,
input [7:0] x1702 ,
input [7:0] x1703 ,
input [7:0] x1704 ,
input [7:0] x1705 ,
input [7:0] x1706 ,
input [7:0] x1707 ,
input [7:0] x1708 ,
input [7:0] x1709 ,
input [7:0] x1710 ,
input [7:0] x1711 ,
input [7:0] x1712 ,
input [7:0] x1713 ,
input [7:0] x1714 ,
input [7:0] x1715 ,
input [7:0] x1716 ,
input [7:0] x1717 ,
input [7:0] x1718 ,
input [7:0] x1719 ,
input [7:0] x1720 ,
input [7:0] x1721 ,
input [7:0] x1722 ,
input [7:0] x1723 ,
input [7:0] x1724 ,
input [7:0] x1725 ,
input [7:0] x1726 ,
input [7:0] x1727 ,
input [7:0] x1728 ,
input [7:0] x1729 ,
input [7:0] x1730 ,
input [7:0] x1731 ,
input [7:0] x1732 ,
input [7:0] x1733 ,
input [7:0] x1734 ,
input [7:0] x1735 ,
input [7:0] x1736 ,
input [7:0] x1737 ,
input [7:0] x1738 ,
input [7:0] x1739 ,
input [7:0] x1740 ,
input [7:0] x1741 ,
input [7:0] x1742 ,
input [7:0] x1743 ,
input [7:0] x1744 ,
input [7:0] x1745 ,
input [7:0] x1746 ,
input [7:0] x1747 ,
input [7:0] x1748 ,
input [7:0] x1749 ,
input [7:0] x1750 ,
input [7:0] x1751 ,
input [7:0] x1752 ,
input [7:0] x1753 ,
input [7:0] x1754 ,
input [7:0] x1755 ,
input [7:0] x1756 ,
input [7:0] x1757 ,
input [7:0] x1758 ,
input [7:0] x1759 ,
input [7:0] x1760 ,
input [7:0] x1761 ,
input [7:0] x1762 ,
input [7:0] x1763 ,
input [7:0] x1764 ,
input [7:0] x1765 ,
input [7:0] x1766 ,
input [7:0] x1767 ,
input [7:0] x1768 ,
input [7:0] x1769 ,
input [7:0] x1770 ,
input [7:0] x1771 ,
input [7:0] x1772 ,
input [7:0] x1773 ,
input [7:0] x1774 ,
input [7:0] x1775 ,
input [7:0] x1776 ,
input [7:0] x1777 ,
input [7:0] x1778 ,
input [7:0] x1779 ,
input [7:0] x1780 ,
input [7:0] x1781 ,
input [7:0] x1782 ,
input [7:0] x1783 ,
input [7:0] x1784 ,
input [7:0] x1785 ,
input [7:0] x1786 ,
input [7:0] x1787 ,
input [7:0] x1788 ,
input [7:0] x1789 ,
input [7:0] x1790 ,
input [7:0] x1791 ,
input [7:0] x1792 ,
input [7:0] x1793 ,
input [7:0] x1794 ,
input [7:0] x1795 ,
input [7:0] x1796 ,
input [7:0] x1797 ,
input [7:0] x1798 ,
input [7:0] x1799 ,
input [7:0] x1800 ,
input [7:0] x1801 ,
input [7:0] x1802 ,
input [7:0] x1803 ,
input [7:0] x1804 ,
input [7:0] x1805 ,
input [7:0] x1806 ,
input [7:0] x1807 ,
input [7:0] x1808 ,
input [7:0] x1809 ,
input [7:0] x1810 ,
input [7:0] x1811 ,
input [7:0] x1812 ,
input [7:0] x1813 ,
input [7:0] x1814 ,
input [7:0] x1815 ,
input [7:0] x1816 ,
input [7:0] x1817 ,
input [7:0] x1818 ,
input [7:0] x1819 ,
input [7:0] x1820 ,
input [7:0] x1821 ,
input [7:0] x1822 ,
input [7:0] x1823 ,
input [7:0] x1824 ,
input [7:0] x1825 ,
input [7:0] x1826 ,
input [7:0] x1827 ,
input [7:0] x1828 ,
input [7:0] x1829 ,
input [7:0] x1830 ,
input [7:0] x1831 ,
input [7:0] x1832 ,
input [7:0] x1833 ,
input [7:0] x1834 ,
input [7:0] x1835 ,
input [7:0] x1836 ,
input [7:0] x1837 ,
input [7:0] x1838 ,
input [7:0] x1839 ,
input [7:0] x1840 ,
input [7:0] x1841 ,
input [7:0] x1842 ,
input [7:0] x1843 ,
input [7:0] x1844 ,
input [7:0] x1845 ,
input [7:0] x1846 ,
input [7:0] x1847 ,
input [7:0] x1848 ,
input [7:0] x1849 ,
input [7:0] x1850 ,
input [7:0] x1851 ,
input [7:0] x1852 ,
input [7:0] x1853 ,
input [7:0] x1854 ,
input [7:0] x1855 ,
input [7:0] x1856 ,
input [7:0] x1857 ,
input [7:0] x1858 ,
input [7:0] x1859 ,
input [7:0] x1860 ,
input [7:0] x1861 ,
input [7:0] x1862 ,
input [7:0] x1863 ,
input [7:0] x1864 ,
input [7:0] x1865 ,
input [7:0] x1866 ,
input [7:0] x1867 ,
input [7:0] x1868 ,
input [7:0] x1869 ,
input [7:0] x1870 ,
input [7:0] x1871 ,
input [7:0] x1872 ,
input [7:0] x1873 ,
input [7:0] x1874 ,
input [7:0] x1875 ,
input [7:0] x1876 ,
input [7:0] x1877 ,
input [7:0] x1878 ,
input [7:0] x1879 ,
input [7:0] x1880 ,
input [7:0] x1881 ,
input [7:0] x1882 ,
input [7:0] x1883 ,
input [7:0] x1884 ,
input [7:0] x1885 ,
input [7:0] x1886 ,
input [7:0] x1887 ,
input [7:0] x1888 ,
input [7:0] x1889 ,
input [7:0] x1890 ,
input [7:0] x1891 ,
input [7:0] x1892 ,
input [7:0] x1893 ,
input [7:0] x1894 ,
input [7:0] x1895 ,
input [7:0] x1896 ,
input [7:0] x1897 ,
input [7:0] x1898 ,
input [7:0] x1899 ,
input [7:0] x1900 ,
input [7:0] x1901 ,
input [7:0] x1902 ,
input [7:0] x1903 ,
input [7:0] x1904 ,
input [7:0] x1905 ,
input [7:0] x1906 ,
input [7:0] x1907 ,
input [7:0] x1908 ,
input [7:0] x1909 ,
input [7:0] x1910 ,
input [7:0] x1911 ,
input [7:0] x1912 ,
input [7:0] x1913 ,
input [7:0] x1914 ,
input [7:0] x1915 ,
input [7:0] x1916 ,
input [7:0] x1917 ,
input [7:0] x1918 ,
input [7:0] x1919 ,
input [7:0] x1920 ,
input [7:0] x1921 ,
input [7:0] x1922 ,
input [7:0] x1923 ,
input [7:0] x1924 ,
input [7:0] x1925 ,
input [7:0] x1926 ,
input [7:0] x1927 ,
input [7:0] x1928 ,
input [7:0] x1929 ,
input [7:0] x1930 ,
input [7:0] x1931 ,
input [7:0] x1932 ,
input [7:0] x1933 ,
input [7:0] x1934 ,
input [7:0] x1935 ,
input [7:0] x1936 ,
input [7:0] x1937 ,
input [7:0] x1938 ,
input [7:0] x1939 ,
input [7:0] x1940 ,
input [7:0] x1941 ,
input [7:0] x1942 ,
input [7:0] x1943 ,
input [7:0] x1944 ,
input [7:0] x1945 ,
input [7:0] x1946 ,
input [7:0] x1947 ,
input [7:0] x1948 ,
input [7:0] x1949 ,
input [7:0] x1950 ,
input [7:0] x1951 ,
input [7:0] x1952 ,
input [7:0] x1953 ,
input [7:0] x1954 ,
input [7:0] x1955 ,
input [7:0] x1956 ,
input [7:0] x1957 ,
input [7:0] x1958 ,
input [7:0] x1959 ,
input [7:0] x1960 ,
input [7:0] x1961 ,
input [7:0] x1962 ,
input [7:0] x1963 ,
input [7:0] x1964 ,
input [7:0] x1965 ,
input [7:0] x1966 ,
input [7:0] x1967 ,
input [7:0] x1968 ,
input [7:0] x1969 ,
input [7:0] x1970 ,
input [7:0] x1971 ,
input [7:0] x1972 ,
input [7:0] x1973 ,
input [7:0] x1974 ,
input [7:0] x1975 ,
input [7:0] x1976 ,
input [7:0] x1977 ,
input [7:0] x1978 ,
input [7:0] x1979 ,
input [7:0] x1980 ,
input [7:0] x1981 ,
input [7:0] x1982 ,
input [7:0] x1983 ,
input [7:0] x1984 ,
input [7:0] x1985 ,
input [7:0] x1986 ,
input [7:0] x1987 ,
input [7:0] x1988 ,
input [7:0] x1989 ,
input [7:0] x1990 ,
input [7:0] x1991 ,
input [7:0] x1992 ,
input [7:0] x1993 ,
input [7:0] x1994 ,
input [7:0] x1995 ,
input [7:0] x1996 ,
input [7:0] x1997 ,
input [7:0] x1998 ,
input [7:0] x1999 ,
input [7:0] x2000 ,
input [7:0] x2001 ,
input [7:0] x2002 ,
input [7:0] x2003 ,
input [7:0] x2004 ,
input [7:0] x2005 ,
input [7:0] x2006 ,
input [7:0] x2007 ,
input [7:0] x2008 ,
input [7:0] x2009 ,
input [7:0] x2010 ,
input [7:0] x2011 ,
input [7:0] x2012 ,
input [7:0] x2013 ,
input [7:0] x2014 ,
input [7:0] x2015 ,
input [7:0] x2016 ,
input [7:0] x2017 ,
input [7:0] x2018 ,
input [7:0] x2019 ,
input [7:0] x2020 ,
input [7:0] x2021 ,
input [7:0] x2022 ,
input [7:0] x2023 ,
input [7:0] x2024 ,
input [7:0] x2025 ,
input [7:0] x2026 ,
input [7:0] x2027 ,
input [7:0] x2028 ,
input [7:0] x2029 ,
input [7:0] x2030 ,
input [7:0] x2031 ,
input [7:0] x2032 ,
input [7:0] x2033 ,
input [7:0] x2034 ,
input [7:0] x2035 ,
input [7:0] x2036 ,
input [7:0] x2037 ,
input [7:0] x2038 ,
input [7:0] x2039 ,
input [7:0] x2040 ,
input [7:0] x2041 ,
input [7:0] x2042 ,
input [7:0] x2043 ,
input [7:0] x2044 ,
input [7:0] x2045 ,
input [7:0] x2046 ,
input [7:0] x2047 ,
input [7:0] x2048 ,
input [7:0] x2049 ,
input [7:0] x2050 ,
input [7:0] x2051 ,
input [7:0] x2052 ,
input [7:0] x2053 ,
input [7:0] x2054 ,
input [7:0] x2055 ,
input [7:0] x2056 ,
input [7:0] x2057 ,
input [7:0] x2058 ,
input [7:0] x2059 ,
input [7:0] x2060 ,
input [7:0] x2061 ,
input [7:0] x2062 ,
input [7:0] x2063 ,
input [7:0] x2064 ,
input [7:0] x2065 ,
input [7:0] x2066 ,
input [7:0] x2067 ,
input [7:0] x2068 ,
input [7:0] x2069 ,
input [7:0] x2070 ,
input [7:0] x2071 ,
input [7:0] x2072 ,
input [7:0] x2073 ,
input [7:0] x2074 ,
input [7:0] x2075 ,
input [7:0] x2076 ,
input [7:0] x2077 ,
input [7:0] x2078 ,
input [7:0] x2079 ,
input [7:0] x2080 ,
input [7:0] x2081 ,
input [7:0] x2082 ,
input [7:0] x2083 ,
input [7:0] x2084 ,
input [7:0] x2085 ,
input [7:0] x2086 ,
input [7:0] x2087 ,
input [7:0] x2088 ,
input [7:0] x2089 ,
input [7:0] x2090 ,
input [7:0] x2091 ,
input [7:0] x2092 ,
input [7:0] x2093 ,
input [7:0] x2094 ,
input [7:0] x2095 ,
input [7:0] x2096 ,
input [7:0] x2097 ,
input [7:0] x2098 ,
input [7:0] x2099 ,
input [7:0] x2100 ,
input [7:0] x2101 ,
input [7:0] x2102 ,
input [7:0] x2103 ,
input [7:0] x2104 ,
input [7:0] x2105 ,
input [7:0] x2106 ,
input [7:0] x2107 ,
input [7:0] x2108 ,
input [7:0] x2109 ,
input [7:0] x2110 ,
input [7:0] x2111 ,
input [7:0] x2112 ,
input [7:0] x2113 ,
input [7:0] x2114 ,
input [7:0] x2115 ,
input [7:0] x2116 ,
input [7:0] x2117 ,
input [7:0] x2118 ,
input [7:0] x2119 ,
input [7:0] x2120 ,
input [7:0] x2121 ,
input [7:0] x2122 ,
input [7:0] x2123 ,
input [7:0] x2124 ,
input [7:0] x2125 ,
input [7:0] x2126 ,
input [7:0] x2127 ,
input [7:0] x2128 ,
input [7:0] x2129 ,
input [7:0] x2130 ,
input [7:0] x2131 ,
input [7:0] x2132 ,
input [7:0] x2133 ,
input [7:0] x2134 ,
input [7:0] x2135 ,
input [7:0] x2136 ,
input [7:0] x2137 ,
input [7:0] x2138 ,
input [7:0] x2139 ,
input [7:0] x2140 ,
input [7:0] x2141 ,
input [7:0] x2142 ,
input [7:0] x2143 ,
input [7:0] x2144 ,
input [7:0] x2145 ,
input [7:0] x2146 ,
input [7:0] x2147 ,
input [7:0] x2148 ,
input [7:0] x2149 ,
input [7:0] x2150 ,
input [7:0] x2151 ,
input [7:0] x2152 ,
input [7:0] x2153 ,
input [7:0] x2154 ,
input [7:0] x2155 ,
input [7:0] x2156 ,
input [7:0] x2157 ,
input [7:0] x2158 ,
input [7:0] x2159 ,
input [7:0] x2160 ,
input [7:0] x2161 ,
input [7:0] x2162 ,
input [7:0] x2163 ,
input [7:0] x2164 ,
input [7:0] x2165 ,
input [7:0] x2166 ,
input [7:0] x2167 ,
input [7:0] x2168 ,
input [7:0] x2169 ,
input [7:0] x2170 ,
input [7:0] x2171 ,
input [7:0] x2172 ,
input [7:0] x2173 ,
input [7:0] x2174 ,
input [7:0] x2175 ,
input [7:0] x2176 ,
input [7:0] x2177 ,
input [7:0] x2178 ,
input [7:0] x2179 ,
input [7:0] x2180 ,
input [7:0] x2181 ,
input [7:0] x2182 ,
input [7:0] x2183 ,
input [7:0] x2184 ,
input [7:0] x2185 ,
input [7:0] x2186 ,
input [7:0] x2187 ,
input [7:0] x2188 ,
input [7:0] x2189 ,
input [7:0] x2190 ,
input [7:0] x2191 ,
input [7:0] x2192 ,
input [7:0] x2193 ,
input [7:0] x2194 ,
input [7:0] x2195 ,
input [7:0] x2196 ,
input [7:0] x2197 ,
input [7:0] x2198 ,
input [7:0] x2199 ,
input [7:0] x2200 ,
input [7:0] x2201 ,
input [7:0] x2202 ,
input [7:0] x2203 ,
input [7:0] x2204 ,
input [7:0] x2205 ,
input [7:0] x2206 ,
input [7:0] x2207 ,
input [7:0] x2208 ,
input [7:0] x2209 ,
input [7:0] x2210 ,
input [7:0] x2211 ,
input [7:0] x2212 ,
input [7:0] x2213 ,
input [7:0] x2214 ,
input [7:0] x2215 ,
input [7:0] x2216 ,
input [7:0] x2217 ,
input [7:0] x2218 ,
input [7:0] x2219 ,
input [7:0] x2220 ,
input [7:0] x2221 ,
input [7:0] x2222 ,
input [7:0] x2223 ,
input [7:0] x2224 ,
input [7:0] x2225 ,
input [7:0] x2226 ,
input [7:0] x2227 ,
input [7:0] x2228 ,
input [7:0] x2229 ,
input [7:0] x2230 ,
input [7:0] x2231 ,
input [7:0] x2232 ,
input [7:0] x2233 ,
input [7:0] x2234 ,
input [7:0] x2235 ,
input [7:0] x2236 ,
input [7:0] x2237 ,
input [7:0] x2238 ,
input [7:0] x2239 ,
input [7:0] x2240 ,
input [7:0] x2241 ,
input [7:0] x2242 ,
input [7:0] x2243 ,
input [7:0] x2244 ,
input [7:0] x2245 ,
input [7:0] x2246 ,
input [7:0] x2247 ,
input [7:0] x2248 ,
input [7:0] x2249 ,
input [7:0] x2250 ,
input [7:0] x2251 ,
input [7:0] x2252 ,
input [7:0] x2253 ,
input [7:0] x2254 ,
input [7:0] x2255 ,
input [7:0] x2256 ,
input [7:0] x2257 ,
input [7:0] x2258 ,
input [7:0] x2259 ,
input [7:0] x2260 ,
input [7:0] x2261 ,
input [7:0] x2262 ,
input [7:0] x2263 ,
input [7:0] x2264 ,
input [7:0] x2265 ,
input [7:0] x2266 ,
input [7:0] x2267 ,
input [7:0] x2268 ,
input [7:0] x2269 ,
input [7:0] x2270 ,
input [7:0] x2271 ,
input [7:0] x2272 ,
input [7:0] x2273 ,
input [7:0] x2274 ,
input [7:0] x2275 ,
input [7:0] x2276 ,
input [7:0] x2277 ,
input [7:0] x2278 ,
input [7:0] x2279 ,
input [7:0] x2280 ,
input [7:0] x2281 ,
input [7:0] x2282 ,
input [7:0] x2283 ,
input [7:0] x2284 ,
input [7:0] x2285 ,
input [7:0] x2286 ,
input [7:0] x2287 ,
input [7:0] x2288 ,
input [7:0] x2289 ,
input [7:0] x2290 ,
input [7:0] x2291 ,
input [7:0] x2292 ,
input [7:0] x2293 ,
input [7:0] x2294 ,
input [7:0] x2295 ,
input [7:0] x2296 ,
input [7:0] x2297 ,
input [7:0] x2298 ,
input [7:0] x2299 ,
input [7:0] x2300 ,
input [7:0] x2301 ,
input [7:0] x2302 ,
input [7:0] x2303 ,
input [7:0] x2304 ,
input [7:0] x2305 ,
input [7:0] x2306 ,
input [7:0] x2307 ,
input [7:0] x2308 ,
input [7:0] x2309 ,
input [7:0] x2310 ,
input [7:0] x2311 ,
input [7:0] x2312 ,
input [7:0] x2313 ,
input [7:0] x2314 ,
input [7:0] x2315 ,
input [7:0] x2316 ,
input [7:0] x2317 ,
input [7:0] x2318 ,
input [7:0] x2319 ,
input [7:0] x2320 ,
input [7:0] x2321 ,
input [7:0] x2322 ,
input [7:0] x2323 ,
input [7:0] x2324 ,
input [7:0] x2325 ,
input [7:0] x2326 ,
input [7:0] x2327 ,
input [7:0] x2328 ,
input [7:0] x2329 ,
input [7:0] x2330 ,
input [7:0] x2331 ,
input [7:0] x2332 ,
input [7:0] x2333 ,
input [7:0] x2334 ,
input [7:0] x2335 ,
input [7:0] x2336 ,
input [7:0] x2337 ,
input [7:0] x2338 ,
input [7:0] x2339 ,
input [7:0] x2340 ,
input [7:0] x2341 ,
input [7:0] x2342 ,
input [7:0] x2343 ,
input [7:0] x2344 ,
input [7:0] x2345 ,
input [7:0] x2346 ,
input [7:0] x2347 ,
input [7:0] x2348 ,
input [7:0] x2349 ,
input [7:0] x2350 ,
input [7:0] x2351 ,
input [7:0] x2352 ,
input [7:0] x2353 ,
input [7:0] x2354 ,
input [7:0] x2355 ,
input [7:0] x2356 ,
input [7:0] x2357 ,
input [7:0] x2358 ,
input [7:0] x2359 ,
input [7:0] x2360 ,
input [7:0] x2361 ,
input [7:0] x2362 ,
input [7:0] x2363 ,
input [7:0] x2364 ,
input [7:0] x2365 ,
input [7:0] x2366 ,
input [7:0] x2367 ,
input [7:0] x2368 ,
input [7:0] x2369 ,
input [7:0] x2370 ,
input [7:0] x2371 ,
input [7:0] x2372 ,
input [7:0] x2373 ,
input [7:0] x2374 ,
input [7:0] x2375 ,
input [7:0] x2376 ,
input [7:0] x2377 ,
input [7:0] x2378 ,
input [7:0] x2379 ,
input [7:0] x2380 ,
input [7:0] x2381 ,
input [7:0] x2382 ,
input [7:0] x2383 ,
input [7:0] x2384 ,
input [7:0] x2385 ,
input [7:0] x2386 ,
input [7:0] x2387 ,
input [7:0] x2388 ,
input [7:0] x2389 ,
input [7:0] x2390 ,
input [7:0] x2391 ,
input [7:0] x2392 ,
input [7:0] x2393 ,
input [7:0] x2394 ,
input [7:0] x2395 ,
input [7:0] x2396 ,
input [7:0] x2397 ,
input [7:0] x2398 ,
input [7:0] x2399 ,
input [7:0] x2400 ,
input [7:0] x2401 ,
input [7:0] x2402 ,
input [7:0] x2403 ,
input [7:0] x2404 ,
input [7:0] x2405 ,
input [7:0] x2406 ,
input [7:0] x2407 ,
input [7:0] x2408 ,
input [7:0] x2409 ,
input [7:0] x2410 ,
input [7:0] x2411 ,
input [7:0] x2412 ,
input [7:0] x2413 ,
input [7:0] x2414 ,
input [7:0] x2415 ,
input [7:0] x2416 ,
input [7:0] x2417 ,
input [7:0] x2418 ,
input [7:0] x2419 ,
input [7:0] x2420 ,
input [7:0] x2421 ,
input [7:0] x2422 ,
input [7:0] x2423 ,
input [7:0] x2424 ,
input [7:0] x2425 ,
input [7:0] x2426 ,
input [7:0] x2427 ,
input [7:0] x2428 ,
input [7:0] x2429 ,
input [7:0] x2430 ,
input [7:0] x2431 ,
input [7:0] x2432 ,
input [7:0] x2433 ,
input [7:0] x2434 ,
input [7:0] x2435 ,
input [7:0] x2436 ,
input [7:0] x2437 ,
input [7:0] x2438 ,
input [7:0] x2439 ,
input [7:0] x2440 ,
input [7:0] x2441 ,
input [7:0] x2442 ,
input [7:0] x2443 ,
input [7:0] x2444 ,
input [7:0] x2445 ,
input [7:0] x2446 ,
input [7:0] x2447 ,
input [7:0] x2448 ,
input [7:0] x2449 ,
input [7:0] x2450 ,
input [7:0] x2451 ,
input [7:0] x2452 ,
input [7:0] x2453 ,
input [7:0] x2454 ,
input [7:0] x2455 ,
input [7:0] x2456 ,
input [7:0] x2457 ,
input [7:0] x2458 ,
input [7:0] x2459 ,
input [7:0] x2460 ,
input [7:0] x2461 ,
input [7:0] x2462 ,
input [7:0] x2463 ,
input [7:0] x2464 ,
input [7:0] x2465 ,
input [7:0] x2466 ,
input [7:0] x2467 ,
input [7:0] x2468 ,
input [7:0] x2469 ,
input [7:0] x2470 ,
input [7:0] x2471 ,
input [7:0] x2472 ,
input [7:0] x2473 ,
input [7:0] x2474 ,
input [7:0] x2475 ,
input [7:0] x2476 ,
input [7:0] x2477 ,
input [7:0] x2478 ,
input [7:0] x2479 ,
input [7:0] x2480 ,
input [7:0] x2481 ,
input [7:0] x2482 ,
input [7:0] x2483 ,
input [7:0] x2484 ,
input [7:0] x2485 ,
input [7:0] x2486 ,
input [7:0] x2487 ,
input [7:0] x2488 ,
input [7:0] x2489 ,
input [7:0] x2490 ,
input [7:0] x2491 ,
input [7:0] x2492 ,
input [7:0] x2493 ,
input [7:0] x2494 ,
input [7:0] x2495 ,
input [7:0] x2496 ,
input [7:0] x2497 ,
input [7:0] x2498 ,
input [7:0] x2499 ,
input [7:0] x2500 ,
input [7:0] x2501 ,
input [7:0] x2502 ,
input [7:0] x2503 ,
input [7:0] x2504 ,
input [7:0] x2505 ,
input [7:0] x2506 ,
input [7:0] x2507 ,
input [7:0] x2508 ,
input [7:0] x2509 ,
input [7:0] x2510 ,
input [7:0] x2511 ,
input [7:0] x2512 ,
input [7:0] x2513 ,
input [7:0] x2514 ,
input [7:0] x2515 ,
input [7:0] x2516 ,
input [7:0] x2517 ,
input [7:0] x2518 ,
input [7:0] x2519 ,
input [7:0] x2520 ,
input [7:0] x2521 ,
input [7:0] x2522 ,
input [7:0] x2523 ,
input [7:0] x2524 ,
input [7:0] x2525 ,
input [7:0] x2526 ,
input [7:0] x2527 ,
input [7:0] x2528 ,
input [7:0] x2529 ,
input [7:0] x2530 ,
input [7:0] x2531 ,
input [7:0] x2532 ,
input [7:0] x2533 ,
input [7:0] x2534 ,
input [7:0] x2535 ,
input [7:0] x2536 ,
input [7:0] x2537 ,
input [7:0] x2538 ,
input [7:0] x2539 ,
input [7:0] x2540 ,
input [7:0] x2541 ,
input [7:0] x2542 ,
input [7:0] x2543 ,
input [7:0] x2544 ,
input [7:0] x2545 ,
input [7:0] x2546 ,
input [7:0] x2547 ,
input [7:0] x2548 ,
input [7:0] x2549 ,
input [7:0] x2550 ,
input [7:0] x2551 ,
input [7:0] x2552 ,
input [7:0] x2553 ,
input [7:0] x2554 ,
input [7:0] x2555 ,
input [7:0] x2556 ,
input [7:0] x2557 ,
input [7:0] x2558 ,
input [7:0] x2559 ,
input [7:0] x2560 ,
input [7:0] x2561 ,
input [7:0] x2562 ,
input [7:0] x2563 ,
input [7:0] x2564 ,
input [7:0] x2565 ,
input [7:0] x2566 ,
input [7:0] x2567 ,
input [7:0] x2568 ,
input [7:0] x2569 ,
input [7:0] x2570 ,
input [7:0] x2571 ,
input [7:0] x2572 ,
input [7:0] x2573 ,
input [7:0] x2574 ,
input [7:0] x2575 ,
input [7:0] x2576 ,
input [7:0] x2577 ,
input [7:0] x2578 ,
input [7:0] x2579 ,
input [7:0] x2580 ,
input [7:0] x2581 ,
input [7:0] x2582 ,
input [7:0] x2583 ,
input [7:0] x2584 ,
input [7:0] x2585 ,
input [7:0] x2586 ,
input [7:0] x2587 ,
input [7:0] x2588 ,
input [7:0] x2589 ,
input [7:0] x2590 ,
input [7:0] x2591 ,
input [7:0] x2592 ,
input [7:0] x2593 ,
input [7:0] x2594 ,
input [7:0] x2595 ,
input [7:0] x2596 ,
input [7:0] x2597 ,
input [7:0] x2598 ,
input [7:0] x2599 ,
input [7:0] x2600 ,
input [7:0] x2601 ,
input [7:0] x2602 ,
input [7:0] x2603 ,
input [7:0] x2604 ,
input [7:0] x2605 ,
input [7:0] x2606 ,
input [7:0] x2607 ,
input [7:0] x2608 ,
input [7:0] x2609 ,
input [7:0] x2610 ,
input [7:0] x2611 ,
input [7:0] x2612 ,
input [7:0] x2613 ,
input [7:0] x2614 ,
input [7:0] x2615 ,
input [7:0] x2616 ,
input [7:0] x2617 ,
input [7:0] x2618 ,
input [7:0] x2619 ,
input [7:0] x2620 ,
input [7:0] x2621 ,
input [7:0] x2622 ,
input [7:0] x2623 ,
input [7:0] x2624 ,
input [7:0] x2625 ,
input [7:0] x2626 ,
input [7:0] x2627 ,
input [7:0] x2628 ,
input [7:0] x2629 ,
input [7:0] x2630 ,
input [7:0] x2631 ,
input [7:0] x2632 ,
input [7:0] x2633 ,
input [7:0] x2634 ,
input [7:0] x2635 ,
input [7:0] x2636 ,
input [7:0] x2637 ,
input [7:0] x2638 ,
input [7:0] x2639 ,
input [7:0] x2640 ,
input [7:0] x2641 ,
input [7:0] x2642 ,
input [7:0] x2643 ,
input [7:0] x2644 ,
input [7:0] x2645 ,
input [7:0] x2646 ,
input [7:0] x2647 ,
input [7:0] x2648 ,
input [7:0] x2649 ,
input [7:0] x2650 ,
input [7:0] x2651 ,
input [7:0] x2652 ,
input [7:0] x2653 ,
input [7:0] x2654 ,
input [7:0] x2655 ,
input [7:0] x2656 ,
input [7:0] x2657 ,
input [7:0] x2658 ,
input [7:0] x2659 ,
input [7:0] x2660 ,
input [7:0] x2661 ,
input [7:0] x2662 ,
input [7:0] x2663 ,
input [7:0] x2664 ,
input [7:0] x2665 ,
input [7:0] x2666 ,
input [7:0] x2667 ,
input [7:0] x2668 ,
input [7:0] x2669 ,
input [7:0] x2670 ,
input [7:0] x2671 ,
input [7:0] x2672 ,
input [7:0] x2673 ,
input [7:0] x2674 ,
input [7:0] x2675 ,
input [7:0] x2676 ,
input [7:0] x2677 ,
input [7:0] x2678 ,
input [7:0] x2679 ,
input [7:0] x2680 ,
input [7:0] x2681 ,
input [7:0] x2682 ,
input [7:0] x2683 ,
input [7:0] x2684 ,
input [7:0] x2685 ,
input [7:0] x2686 ,
input [7:0] x2687 ,
input [7:0] x2688 ,
input [7:0] x2689 ,
input [7:0] x2690 ,
input [7:0] x2691 ,
input [7:0] x2692 ,
input [7:0] x2693 ,
input [7:0] x2694 ,
input [7:0] x2695 ,
input [7:0] x2696 ,
input [7:0] x2697 ,
input [7:0] x2698 ,
input [7:0] x2699 ,
input [7:0] x2700 ,
input [7:0] x2701 ,
input [7:0] x2702 ,
input [7:0] x2703 ,
input [7:0] x2704 ,
input [7:0] x2705 ,
input [7:0] x2706 ,
input [7:0] x2707 ,
input [7:0] x2708 ,
input [7:0] x2709 ,
input [7:0] x2710 ,
input [7:0] x2711 ,
input [7:0] x2712 ,
input [7:0] x2713 ,
input [7:0] x2714 ,
input [7:0] x2715 ,
input [7:0] x2716 ,
input [7:0] x2717 ,
input [7:0] x2718 ,
input [7:0] x2719 ,
input [7:0] x2720 ,
input [7:0] x2721 ,
input [7:0] x2722 ,
input [7:0] x2723 ,
input [7:0] x2724 ,
input [7:0] x2725 ,
input [7:0] x2726 ,
input [7:0] x2727 ,
input [7:0] x2728 ,
input [7:0] x2729 ,
input [7:0] x2730 ,
input [7:0] x2731 ,
input [7:0] x2732 ,
input [7:0] x2733 ,
input [7:0] x2734 ,
input [7:0] x2735 ,
input [7:0] x2736 ,
input [7:0] x2737 ,
input [7:0] x2738 ,
input [7:0] x2739 ,
input [7:0] x2740 ,
input [7:0] x2741 ,
input [7:0] x2742 ,
input [7:0] x2743 ,
input [7:0] x2744 ,
input [7:0] x2745 ,
input [7:0] x2746 ,
input [7:0] x2747 ,
input [7:0] x2748 ,
input [7:0] x2749 ,
input [7:0] x2750 ,
input [7:0] x2751 ,
input [7:0] x2752 ,
input [7:0] x2753 ,
input [7:0] x2754 ,
input [7:0] x2755 ,
input [7:0] x2756 ,
input [7:0] x2757 ,
input [7:0] x2758 ,
input [7:0] x2759 ,
input [7:0] x2760 ,
input [7:0] x2761 ,
input [7:0] x2762 ,
input [7:0] x2763 ,
input [7:0] x2764 ,
input [7:0] x2765 ,
input [7:0] x2766 ,
input [7:0] x2767 ,
input [7:0] x2768 ,
input [7:0] x2769 ,
input [7:0] x2770 ,
input [7:0] x2771 ,
input [7:0] x2772 ,
input [7:0] x2773 ,
input [7:0] x2774 ,
input [7:0] x2775 ,
input [7:0] x2776 ,
input [7:0] x2777 ,
input [7:0] x2778 ,
input [7:0] x2779 ,
input [7:0] x2780 ,
input [7:0] x2781 ,
input [7:0] x2782 ,
input [7:0] x2783 ,
input [7:0] x2784 ,
input [7:0] x2785 ,
input [7:0] x2786 ,
input [7:0] x2787 ,
input [7:0] x2788 ,
input [7:0] x2789 ,
input [7:0] x2790 ,
input [7:0] x2791 ,
input [7:0] x2792 ,
input [7:0] x2793 ,
input [7:0] x2794 ,
input [7:0] x2795 ,
input [7:0] x2796 ,
input [7:0] x2797 ,
input [7:0] x2798 ,
input [7:0] x2799 ,
input [7:0] x2800 ,
input [7:0] x2801 ,
input [7:0] x2802 ,
input [7:0] x2803 ,
input [7:0] x2804 ,
input [7:0] x2805 ,
input [7:0] x2806 ,
input [7:0] x2807 ,
input [7:0] x2808 ,
input [7:0] x2809 ,
input [7:0] x2810 ,
input [7:0] x2811 ,
input [7:0] x2812 ,
input [7:0] x2813 ,
input [7:0] x2814 ,
input [7:0] x2815 ,
input [7:0] x2816 ,
input [7:0] x2817 ,
input [7:0] x2818 ,
input [7:0] x2819 ,
input [7:0] x2820 ,
input [7:0] x2821 ,
input [7:0] x2822 ,
input [7:0] x2823 ,
input [7:0] x2824 ,
input [7:0] x2825 ,
input [7:0] x2826 ,
input [7:0] x2827 ,
input [7:0] x2828 ,
input [7:0] x2829 ,
input [7:0] x2830 ,
input [7:0] x2831 ,
input [7:0] x2832 ,
input [7:0] x2833 ,
input [7:0] x2834 ,
input [7:0] x2835 ,
input [7:0] x2836 ,
input [7:0] x2837 ,
input [7:0] x2838 ,
input [7:0] x2839 ,
input [7:0] x2840 ,
input [7:0] x2841 ,
input [7:0] x2842 ,
input [7:0] x2843 ,
input [7:0] x2844 ,
input [7:0] x2845 ,
input [7:0] x2846 ,
input [7:0] x2847 ,
input [7:0] x2848 ,
input [7:0] x2849 ,
input [7:0] x2850 ,
input [7:0] x2851 ,
input [7:0] x2852 ,
input [7:0] x2853 ,
input [7:0] x2854 ,
input [7:0] x2855 ,
input [7:0] x2856 ,
input [7:0] x2857 ,
input [7:0] x2858 ,
input [7:0] x2859 ,
input [7:0] x2860 ,
input [7:0] x2861 ,
input [7:0] x2862 ,
input [7:0] x2863 ,
input [7:0] x2864 ,
input [7:0] x2865 ,
input [7:0] x2866 ,
input [7:0] x2867 ,
input [7:0] x2868 ,
input [7:0] x2869 ,
input [7:0] x2870 ,
input [7:0] x2871 ,
input [7:0] x2872 ,
input [7:0] x2873 ,
input [7:0] x2874 ,
input [7:0] x2875 ,
input [7:0] x2876 ,
input [7:0] x2877 ,
input [7:0] x2878 ,
input [7:0] x2879 ,
input [7:0] x2880 ,
input [7:0] x2881 ,
input [7:0] x2882 ,
input [7:0] x2883 ,
input [7:0] x2884 ,
input [7:0] x2885 ,
input [7:0] x2886 ,
input [7:0] x2887 ,
input [7:0] x2888 ,
input [7:0] x2889 ,
input [7:0] x2890 ,
input [7:0] x2891 ,
input [7:0] x2892 ,
input [7:0] x2893 ,
input [7:0] x2894 ,
input [7:0] x2895 ,
input [7:0] x2896 ,
input [7:0] x2897 ,
input [7:0] x2898 ,
input [7:0] x2899 ,
input [7:0] x2900 ,
input [7:0] x2901 ,
input [7:0] x2902 ,
input [7:0] x2903 ,
input [7:0] x2904 ,
input [7:0] x2905 ,
input [7:0] x2906 ,
input [7:0] x2907 ,
input [7:0] x2908 ,
input [7:0] x2909 ,
input [7:0] x2910 ,
input [7:0] x2911 ,
input [7:0] x2912 ,
input [7:0] x2913 ,
input [7:0] x2914 ,
input [7:0] x2915 ,
input [7:0] x2916 ,
input [7:0] x2917 ,
input [7:0] x2918 ,
input [7:0] x2919 ,
input [7:0] x2920 ,
input [7:0] x2921 ,
input [7:0] x2922 ,
input [7:0] x2923 ,
input [7:0] x2924 ,
input [7:0] x2925 ,
input [7:0] x2926 ,
input [7:0] x2927 ,
input [7:0] x2928 ,
input [7:0] x2929 ,
input [7:0] x2930 ,
input [7:0] x2931 ,
input [7:0] x2932 ,
input [7:0] x2933 ,
input [7:0] x2934 ,
input [7:0] x2935 ,
input [7:0] x2936 ,
input [7:0] x2937 ,
input [7:0] x2938 ,
input [7:0] x2939 ,
input [7:0] x2940 ,
input [7:0] x2941 ,
input [7:0] x2942 ,
input [7:0] x2943 ,
input [7:0] x2944 ,
input [7:0] x2945 ,
input [7:0] x2946 ,
input [7:0] x2947 ,
input [7:0] x2948 ,
input [7:0] x2949 ,
input [7:0] x2950 ,
input [7:0] x2951 ,
input [7:0] x2952 ,
input [7:0] x2953 ,
input [7:0] x2954 ,
input [7:0] x2955 ,
input [7:0] x2956 ,
input [7:0] x2957 ,
input [7:0] x2958 ,
input [7:0] x2959 ,
input [7:0] x2960 ,
input [7:0] x2961 ,
input [7:0] x2962 ,
input [7:0] x2963 ,
input [7:0] x2964 ,
input [7:0] x2965 ,
input [7:0] x2966 ,
input [7:0] x2967 ,
input [7:0] x2968 ,
input [7:0] x2969 ,
input [7:0] x2970 ,
input [7:0] x2971 ,
input [7:0] x2972 ,
input [7:0] x2973 ,
input [7:0] x2974 ,
input [7:0] x2975 ,
input [7:0] x2976 ,
input [7:0] x2977 ,
input [7:0] x2978 ,
input [7:0] x2979 ,
input [7:0] x2980 ,
input [7:0] x2981 ,
input [7:0] x2982 ,
input [7:0] x2983 ,
input [7:0] x2984 ,
input [7:0] x2985 ,
input [7:0] x2986 ,
input [7:0] x2987 ,
input [7:0] x2988 ,
input [7:0] x2989 ,
input [7:0] x2990 ,
input [7:0] x2991 ,
input [7:0] x2992 ,
input [7:0] x2993 ,
input [7:0] x2994 ,
input [7:0] x2995 ,
input [7:0] x2996 ,
input [7:0] x2997 ,
input [7:0] x2998 ,
input [7:0] x2999 ,
input [7:0] x3000 ,
input [7:0] x3001 ,
input [7:0] x3002 ,
input [7:0] x3003 ,
input [7:0] x3004 ,
input [7:0] x3005 ,
input [7:0] x3006 ,
input [7:0] x3007 ,
input [7:0] x3008 ,
input [7:0] x3009 ,
input [7:0] x3010 ,
input [7:0] x3011 ,
input [7:0] x3012 ,
input [7:0] x3013 ,
input [7:0] x3014 ,
input [7:0] x3015 ,
input [7:0] x3016 ,
input [7:0] x3017 ,
input [7:0] x3018 ,
input [7:0] x3019 ,
input [7:0] x3020 ,
input [7:0] x3021 ,
input [7:0] x3022 ,
input [7:0] x3023 ,
input [7:0] x3024 ,
input [7:0] x3025 ,
input [7:0] x3026 ,
input [7:0] x3027 ,
input [7:0] x3028 ,
input [7:0] x3029 ,
input [7:0] x3030 ,
input [7:0] x3031 ,
input [7:0] x3032 ,
input [7:0] x3033 ,
input [7:0] x3034 ,
input [7:0] x3035 ,
input [7:0] x3036 ,
input [7:0] x3037 ,
input [7:0] x3038 ,
input [7:0] x3039 ,
input [7:0] x3040 ,
input [7:0] x3041 ,
input [7:0] x3042 ,
input [7:0] x3043 ,
input [7:0] x3044 ,
input [7:0] x3045 ,
input [7:0] x3046 ,
input [7:0] x3047 ,
input [7:0] x3048 ,
input [7:0] x3049 ,
input [7:0] x3050 ,
input [7:0] x3051 ,
input [7:0] x3052 ,
input [7:0] x3053 ,
input [7:0] x3054 ,
input [7:0] x3055 ,
input [7:0] x3056 ,
input [7:0] x3057 ,
input [7:0] x3058 ,
input [7:0] x3059 ,
input [7:0] x3060 ,
input [7:0] x3061 ,
input [7:0] x3062 ,
input [7:0] x3063 ,
input [7:0] x3064 ,
input [7:0] x3065 ,
input [7:0] x3066 ,
input [7:0] x3067 ,
input [7:0] x3068 ,
input [7:0] x3069 ,
input [7:0] x3070 ,
input [7:0] x3071 ,
output [9:0] y 
);
wire [6:0]conv11in[0:16*16*3-1];
Bind b(.x0(x0),
.x1(x1),
.x2(x2),
.x3(x3),
.x4(x4),
.x5(x5),
.x6(x6),
.x7(x7),
.x8(x8),
.x9(x9),
.x10(x10),
.x11(x11),
.x12(x12),
.x13(x13),
.x14(x14),
.x15(x15),
.x16(x16),
.x17(x17),
.x18(x18),
.x19(x19),
.x20(x20),
.x21(x21),
.x22(x22),
.x23(x23),
.x24(x24),
.x25(x25),
.x26(x26),
.x27(x27),
.x28(x28),
.x29(x29),
.x30(x30),
.x31(x31),
.x32(x32),
.x33(x33),
.x34(x34),
.x35(x35),
.x36(x36),
.x37(x37),
.x38(x38),
.x39(x39),
.x40(x40),
.x41(x41),
.x42(x42),
.x43(x43),
.x44(x44),
.x45(x45),
.x46(x46),
.x47(x47),
.x48(x48),
.x49(x49),
.x50(x50),
.x51(x51),
.x52(x52),
.x53(x53),
.x54(x54),
.x55(x55),
.x56(x56),
.x57(x57),
.x58(x58),
.x59(x59),
.x60(x60),
.x61(x61),
.x62(x62),
.x63(x63),
.x64(x64),
.x65(x65),
.x66(x66),
.x67(x67),
.x68(x68),
.x69(x69),
.x70(x70),
.x71(x71),
.x72(x72),
.x73(x73),
.x74(x74),
.x75(x75),
.x76(x76),
.x77(x77),
.x78(x78),
.x79(x79),
.x80(x80),
.x81(x81),
.x82(x82),
.x83(x83),
.x84(x84),
.x85(x85),
.x86(x86),
.x87(x87),
.x88(x88),
.x89(x89),
.x90(x90),
.x91(x91),
.x92(x92),
.x93(x93),
.x94(x94),
.x95(x95),
.x96(x96),
.x97(x97),
.x98(x98),
.x99(x99),
.x100(x100),
.x101(x101),
.x102(x102),
.x103(x103),
.x104(x104),
.x105(x105),
.x106(x106),
.x107(x107),
.x108(x108),
.x109(x109),
.x110(x110),
.x111(x111),
.x112(x112),
.x113(x113),
.x114(x114),
.x115(x115),
.x116(x116),
.x117(x117),
.x118(x118),
.x119(x119),
.x120(x120),
.x121(x121),
.x122(x122),
.x123(x123),
.x124(x124),
.x125(x125),
.x126(x126),
.x127(x127),
.x128(x128),
.x129(x129),
.x130(x130),
.x131(x131),
.x132(x132),
.x133(x133),
.x134(x134),
.x135(x135),
.x136(x136),
.x137(x137),
.x138(x138),
.x139(x139),
.x140(x140),
.x141(x141),
.x142(x142),
.x143(x143),
.x144(x144),
.x145(x145),
.x146(x146),
.x147(x147),
.x148(x148),
.x149(x149),
.x150(x150),
.x151(x151),
.x152(x152),
.x153(x153),
.x154(x154),
.x155(x155),
.x156(x156),
.x157(x157),
.x158(x158),
.x159(x159),
.x160(x160),
.x161(x161),
.x162(x162),
.x163(x163),
.x164(x164),
.x165(x165),
.x166(x166),
.x167(x167),
.x168(x168),
.x169(x169),
.x170(x170),
.x171(x171),
.x172(x172),
.x173(x173),
.x174(x174),
.x175(x175),
.x176(x176),
.x177(x177),
.x178(x178),
.x179(x179),
.x180(x180),
.x181(x181),
.x182(x182),
.x183(x183),
.x184(x184),
.x185(x185),
.x186(x186),
.x187(x187),
.x188(x188),
.x189(x189),
.x190(x190),
.x191(x191),
.x192(x192),
.x193(x193),
.x194(x194),
.x195(x195),
.x196(x196),
.x197(x197),
.x198(x198),
.x199(x199),
.x200(x200),
.x201(x201),
.x202(x202),
.x203(x203),
.x204(x204),
.x205(x205),
.x206(x206),
.x207(x207),
.x208(x208),
.x209(x209),
.x210(x210),
.x211(x211),
.x212(x212),
.x213(x213),
.x214(x214),
.x215(x215),
.x216(x216),
.x217(x217),
.x218(x218),
.x219(x219),
.x220(x220),
.x221(x221),
.x222(x222),
.x223(x223),
.x224(x224),
.x225(x225),
.x226(x226),
.x227(x227),
.x228(x228),
.x229(x229),
.x230(x230),
.x231(x231),
.x232(x232),
.x233(x233),
.x234(x234),
.x235(x235),
.x236(x236),
.x237(x237),
.x238(x238),
.x239(x239),
.x240(x240),
.x241(x241),
.x242(x242),
.x243(x243),
.x244(x244),
.x245(x245),
.x246(x246),
.x247(x247),
.x248(x248),
.x249(x249),
.x250(x250),
.x251(x251),
.x252(x252),
.x253(x253),
.x254(x254),
.x255(x255),
.x256(x256),
.x257(x257),
.x258(x258),
.x259(x259),
.x260(x260),
.x261(x261),
.x262(x262),
.x263(x263),
.x264(x264),
.x265(x265),
.x266(x266),
.x267(x267),
.x268(x268),
.x269(x269),
.x270(x270),
.x271(x271),
.x272(x272),
.x273(x273),
.x274(x274),
.x275(x275),
.x276(x276),
.x277(x277),
.x278(x278),
.x279(x279),
.x280(x280),
.x281(x281),
.x282(x282),
.x283(x283),
.x284(x284),
.x285(x285),
.x286(x286),
.x287(x287),
.x288(x288),
.x289(x289),
.x290(x290),
.x291(x291),
.x292(x292),
.x293(x293),
.x294(x294),
.x295(x295),
.x296(x296),
.x297(x297),
.x298(x298),
.x299(x299),
.x300(x300),
.x301(x301),
.x302(x302),
.x303(x303),
.x304(x304),
.x305(x305),
.x306(x306),
.x307(x307),
.x308(x308),
.x309(x309),
.x310(x310),
.x311(x311),
.x312(x312),
.x313(x313),
.x314(x314),
.x315(x315),
.x316(x316),
.x317(x317),
.x318(x318),
.x319(x319),
.x320(x320),
.x321(x321),
.x322(x322),
.x323(x323),
.x324(x324),
.x325(x325),
.x326(x326),
.x327(x327),
.x328(x328),
.x329(x329),
.x330(x330),
.x331(x331),
.x332(x332),
.x333(x333),
.x334(x334),
.x335(x335),
.x336(x336),
.x337(x337),
.x338(x338),
.x339(x339),
.x340(x340),
.x341(x341),
.x342(x342),
.x343(x343),
.x344(x344),
.x345(x345),
.x346(x346),
.x347(x347),
.x348(x348),
.x349(x349),
.x350(x350),
.x351(x351),
.x352(x352),
.x353(x353),
.x354(x354),
.x355(x355),
.x356(x356),
.x357(x357),
.x358(x358),
.x359(x359),
.x360(x360),
.x361(x361),
.x362(x362),
.x363(x363),
.x364(x364),
.x365(x365),
.x366(x366),
.x367(x367),
.x368(x368),
.x369(x369),
.x370(x370),
.x371(x371),
.x372(x372),
.x373(x373),
.x374(x374),
.x375(x375),
.x376(x376),
.x377(x377),
.x378(x378),
.x379(x379),
.x380(x380),
.x381(x381),
.x382(x382),
.x383(x383),
.x384(x384),
.x385(x385),
.x386(x386),
.x387(x387),
.x388(x388),
.x389(x389),
.x390(x390),
.x391(x391),
.x392(x392),
.x393(x393),
.x394(x394),
.x395(x395),
.x396(x396),
.x397(x397),
.x398(x398),
.x399(x399),
.x400(x400),
.x401(x401),
.x402(x402),
.x403(x403),
.x404(x404),
.x405(x405),
.x406(x406),
.x407(x407),
.x408(x408),
.x409(x409),
.x410(x410),
.x411(x411),
.x412(x412),
.x413(x413),
.x414(x414),
.x415(x415),
.x416(x416),
.x417(x417),
.x418(x418),
.x419(x419),
.x420(x420),
.x421(x421),
.x422(x422),
.x423(x423),
.x424(x424),
.x425(x425),
.x426(x426),
.x427(x427),
.x428(x428),
.x429(x429),
.x430(x430),
.x431(x431),
.x432(x432),
.x433(x433),
.x434(x434),
.x435(x435),
.x436(x436),
.x437(x437),
.x438(x438),
.x439(x439),
.x440(x440),
.x441(x441),
.x442(x442),
.x443(x443),
.x444(x444),
.x445(x445),
.x446(x446),
.x447(x447),
.x448(x448),
.x449(x449),
.x450(x450),
.x451(x451),
.x452(x452),
.x453(x453),
.x454(x454),
.x455(x455),
.x456(x456),
.x457(x457),
.x458(x458),
.x459(x459),
.x460(x460),
.x461(x461),
.x462(x462),
.x463(x463),
.x464(x464),
.x465(x465),
.x466(x466),
.x467(x467),
.x468(x468),
.x469(x469),
.x470(x470),
.x471(x471),
.x472(x472),
.x473(x473),
.x474(x474),
.x475(x475),
.x476(x476),
.x477(x477),
.x478(x478),
.x479(x479),
.x480(x480),
.x481(x481),
.x482(x482),
.x483(x483),
.x484(x484),
.x485(x485),
.x486(x486),
.x487(x487),
.x488(x488),
.x489(x489),
.x490(x490),
.x491(x491),
.x492(x492),
.x493(x493),
.x494(x494),
.x495(x495),
.x496(x496),
.x497(x497),
.x498(x498),
.x499(x499),
.x500(x500),
.x501(x501),
.x502(x502),
.x503(x503),
.x504(x504),
.x505(x505),
.x506(x506),
.x507(x507),
.x508(x508),
.x509(x509),
.x510(x510),
.x511(x511),
.x512(x512),
.x513(x513),
.x514(x514),
.x515(x515),
.x516(x516),
.x517(x517),
.x518(x518),
.x519(x519),
.x520(x520),
.x521(x521),
.x522(x522),
.x523(x523),
.x524(x524),
.x525(x525),
.x526(x526),
.x527(x527),
.x528(x528),
.x529(x529),
.x530(x530),
.x531(x531),
.x532(x532),
.x533(x533),
.x534(x534),
.x535(x535),
.x536(x536),
.x537(x537),
.x538(x538),
.x539(x539),
.x540(x540),
.x541(x541),
.x542(x542),
.x543(x543),
.x544(x544),
.x545(x545),
.x546(x546),
.x547(x547),
.x548(x548),
.x549(x549),
.x550(x550),
.x551(x551),
.x552(x552),
.x553(x553),
.x554(x554),
.x555(x555),
.x556(x556),
.x557(x557),
.x558(x558),
.x559(x559),
.x560(x560),
.x561(x561),
.x562(x562),
.x563(x563),
.x564(x564),
.x565(x565),
.x566(x566),
.x567(x567),
.x568(x568),
.x569(x569),
.x570(x570),
.x571(x571),
.x572(x572),
.x573(x573),
.x574(x574),
.x575(x575),
.x576(x576),
.x577(x577),
.x578(x578),
.x579(x579),
.x580(x580),
.x581(x581),
.x582(x582),
.x583(x583),
.x584(x584),
.x585(x585),
.x586(x586),
.x587(x587),
.x588(x588),
.x589(x589),
.x590(x590),
.x591(x591),
.x592(x592),
.x593(x593),
.x594(x594),
.x595(x595),
.x596(x596),
.x597(x597),
.x598(x598),
.x599(x599),
.x600(x600),
.x601(x601),
.x602(x602),
.x603(x603),
.x604(x604),
.x605(x605),
.x606(x606),
.x607(x607),
.x608(x608),
.x609(x609),
.x610(x610),
.x611(x611),
.x612(x612),
.x613(x613),
.x614(x614),
.x615(x615),
.x616(x616),
.x617(x617),
.x618(x618),
.x619(x619),
.x620(x620),
.x621(x621),
.x622(x622),
.x623(x623),
.x624(x624),
.x625(x625),
.x626(x626),
.x627(x627),
.x628(x628),
.x629(x629),
.x630(x630),
.x631(x631),
.x632(x632),
.x633(x633),
.x634(x634),
.x635(x635),
.x636(x636),
.x637(x637),
.x638(x638),
.x639(x639),
.x640(x640),
.x641(x641),
.x642(x642),
.x643(x643),
.x644(x644),
.x645(x645),
.x646(x646),
.x647(x647),
.x648(x648),
.x649(x649),
.x650(x650),
.x651(x651),
.x652(x652),
.x653(x653),
.x654(x654),
.x655(x655),
.x656(x656),
.x657(x657),
.x658(x658),
.x659(x659),
.x660(x660),
.x661(x661),
.x662(x662),
.x663(x663),
.x664(x664),
.x665(x665),
.x666(x666),
.x667(x667),
.x668(x668),
.x669(x669),
.x670(x670),
.x671(x671),
.x672(x672),
.x673(x673),
.x674(x674),
.x675(x675),
.x676(x676),
.x677(x677),
.x678(x678),
.x679(x679),
.x680(x680),
.x681(x681),
.x682(x682),
.x683(x683),
.x684(x684),
.x685(x685),
.x686(x686),
.x687(x687),
.x688(x688),
.x689(x689),
.x690(x690),
.x691(x691),
.x692(x692),
.x693(x693),
.x694(x694),
.x695(x695),
.x696(x696),
.x697(x697),
.x698(x698),
.x699(x699),
.x700(x700),
.x701(x701),
.x702(x702),
.x703(x703),
.x704(x704),
.x705(x705),
.x706(x706),
.x707(x707),
.x708(x708),
.x709(x709),
.x710(x710),
.x711(x711),
.x712(x712),
.x713(x713),
.x714(x714),
.x715(x715),
.x716(x716),
.x717(x717),
.x718(x718),
.x719(x719),
.x720(x720),
.x721(x721),
.x722(x722),
.x723(x723),
.x724(x724),
.x725(x725),
.x726(x726),
.x727(x727),
.x728(x728),
.x729(x729),
.x730(x730),
.x731(x731),
.x732(x732),
.x733(x733),
.x734(x734),
.x735(x735),
.x736(x736),
.x737(x737),
.x738(x738),
.x739(x739),
.x740(x740),
.x741(x741),
.x742(x742),
.x743(x743),
.x744(x744),
.x745(x745),
.x746(x746),
.x747(x747),
.x748(x748),
.x749(x749),
.x750(x750),
.x751(x751),
.x752(x752),
.x753(x753),
.x754(x754),
.x755(x755),
.x756(x756),
.x757(x757),
.x758(x758),
.x759(x759),
.x760(x760),
.x761(x761),
.x762(x762),
.x763(x763),
.x764(x764),
.x765(x765),
.x766(x766),
.x767(x767),
.x768(x768),
.x769(x769),
.x770(x770),
.x771(x771),
.x772(x772),
.x773(x773),
.x774(x774),
.x775(x775),
.x776(x776),
.x777(x777),
.x778(x778),
.x779(x779),
.x780(x780),
.x781(x781),
.x782(x782),
.x783(x783),
.x784(x784),
.x785(x785),
.x786(x786),
.x787(x787),
.x788(x788),
.x789(x789),
.x790(x790),
.x791(x791),
.x792(x792),
.x793(x793),
.x794(x794),
.x795(x795),
.x796(x796),
.x797(x797),
.x798(x798),
.x799(x799),
.x800(x800),
.x801(x801),
.x802(x802),
.x803(x803),
.x804(x804),
.x805(x805),
.x806(x806),
.x807(x807),
.x808(x808),
.x809(x809),
.x810(x810),
.x811(x811),
.x812(x812),
.x813(x813),
.x814(x814),
.x815(x815),
.x816(x816),
.x817(x817),
.x818(x818),
.x819(x819),
.x820(x820),
.x821(x821),
.x822(x822),
.x823(x823),
.x824(x824),
.x825(x825),
.x826(x826),
.x827(x827),
.x828(x828),
.x829(x829),
.x830(x830),
.x831(x831),
.x832(x832),
.x833(x833),
.x834(x834),
.x835(x835),
.x836(x836),
.x837(x837),
.x838(x838),
.x839(x839),
.x840(x840),
.x841(x841),
.x842(x842),
.x843(x843),
.x844(x844),
.x845(x845),
.x846(x846),
.x847(x847),
.x848(x848),
.x849(x849),
.x850(x850),
.x851(x851),
.x852(x852),
.x853(x853),
.x854(x854),
.x855(x855),
.x856(x856),
.x857(x857),
.x858(x858),
.x859(x859),
.x860(x860),
.x861(x861),
.x862(x862),
.x863(x863),
.x864(x864),
.x865(x865),
.x866(x866),
.x867(x867),
.x868(x868),
.x869(x869),
.x870(x870),
.x871(x871),
.x872(x872),
.x873(x873),
.x874(x874),
.x875(x875),
.x876(x876),
.x877(x877),
.x878(x878),
.x879(x879),
.x880(x880),
.x881(x881),
.x882(x882),
.x883(x883),
.x884(x884),
.x885(x885),
.x886(x886),
.x887(x887),
.x888(x888),
.x889(x889),
.x890(x890),
.x891(x891),
.x892(x892),
.x893(x893),
.x894(x894),
.x895(x895),
.x896(x896),
.x897(x897),
.x898(x898),
.x899(x899),
.x900(x900),
.x901(x901),
.x902(x902),
.x903(x903),
.x904(x904),
.x905(x905),
.x906(x906),
.x907(x907),
.x908(x908),
.x909(x909),
.x910(x910),
.x911(x911),
.x912(x912),
.x913(x913),
.x914(x914),
.x915(x915),
.x916(x916),
.x917(x917),
.x918(x918),
.x919(x919),
.x920(x920),
.x921(x921),
.x922(x922),
.x923(x923),
.x924(x924),
.x925(x925),
.x926(x926),
.x927(x927),
.x928(x928),
.x929(x929),
.x930(x930),
.x931(x931),
.x932(x932),
.x933(x933),
.x934(x934),
.x935(x935),
.x936(x936),
.x937(x937),
.x938(x938),
.x939(x939),
.x940(x940),
.x941(x941),
.x942(x942),
.x943(x943),
.x944(x944),
.x945(x945),
.x946(x946),
.x947(x947),
.x948(x948),
.x949(x949),
.x950(x950),
.x951(x951),
.x952(x952),
.x953(x953),
.x954(x954),
.x955(x955),
.x956(x956),
.x957(x957),
.x958(x958),
.x959(x959),
.x960(x960),
.x961(x961),
.x962(x962),
.x963(x963),
.x964(x964),
.x965(x965),
.x966(x966),
.x967(x967),
.x968(x968),
.x969(x969),
.x970(x970),
.x971(x971),
.x972(x972),
.x973(x973),
.x974(x974),
.x975(x975),
.x976(x976),
.x977(x977),
.x978(x978),
.x979(x979),
.x980(x980),
.x981(x981),
.x982(x982),
.x983(x983),
.x984(x984),
.x985(x985),
.x986(x986),
.x987(x987),
.x988(x988),
.x989(x989),
.x990(x990),
.x991(x991),
.x992(x992),
.x993(x993),
.x994(x994),
.x995(x995),
.x996(x996),
.x997(x997),
.x998(x998),
.x999(x999),
.x1000(x1000),
.x1001(x1001),
.x1002(x1002),
.x1003(x1003),
.x1004(x1004),
.x1005(x1005),
.x1006(x1006),
.x1007(x1007),
.x1008(x1008),
.x1009(x1009),
.x1010(x1010),
.x1011(x1011),
.x1012(x1012),
.x1013(x1013),
.x1014(x1014),
.x1015(x1015),
.x1016(x1016),
.x1017(x1017),
.x1018(x1018),
.x1019(x1019),
.x1020(x1020),
.x1021(x1021),
.x1022(x1022),
.x1023(x1023),
.x1024(x1024),
.x1025(x1025),
.x1026(x1026),
.x1027(x1027),
.x1028(x1028),
.x1029(x1029),
.x1030(x1030),
.x1031(x1031),
.x1032(x1032),
.x1033(x1033),
.x1034(x1034),
.x1035(x1035),
.x1036(x1036),
.x1037(x1037),
.x1038(x1038),
.x1039(x1039),
.x1040(x1040),
.x1041(x1041),
.x1042(x1042),
.x1043(x1043),
.x1044(x1044),
.x1045(x1045),
.x1046(x1046),
.x1047(x1047),
.x1048(x1048),
.x1049(x1049),
.x1050(x1050),
.x1051(x1051),
.x1052(x1052),
.x1053(x1053),
.x1054(x1054),
.x1055(x1055),
.x1056(x1056),
.x1057(x1057),
.x1058(x1058),
.x1059(x1059),
.x1060(x1060),
.x1061(x1061),
.x1062(x1062),
.x1063(x1063),
.x1064(x1064),
.x1065(x1065),
.x1066(x1066),
.x1067(x1067),
.x1068(x1068),
.x1069(x1069),
.x1070(x1070),
.x1071(x1071),
.x1072(x1072),
.x1073(x1073),
.x1074(x1074),
.x1075(x1075),
.x1076(x1076),
.x1077(x1077),
.x1078(x1078),
.x1079(x1079),
.x1080(x1080),
.x1081(x1081),
.x1082(x1082),
.x1083(x1083),
.x1084(x1084),
.x1085(x1085),
.x1086(x1086),
.x1087(x1087),
.x1088(x1088),
.x1089(x1089),
.x1090(x1090),
.x1091(x1091),
.x1092(x1092),
.x1093(x1093),
.x1094(x1094),
.x1095(x1095),
.x1096(x1096),
.x1097(x1097),
.x1098(x1098),
.x1099(x1099),
.x1100(x1100),
.x1101(x1101),
.x1102(x1102),
.x1103(x1103),
.x1104(x1104),
.x1105(x1105),
.x1106(x1106),
.x1107(x1107),
.x1108(x1108),
.x1109(x1109),
.x1110(x1110),
.x1111(x1111),
.x1112(x1112),
.x1113(x1113),
.x1114(x1114),
.x1115(x1115),
.x1116(x1116),
.x1117(x1117),
.x1118(x1118),
.x1119(x1119),
.x1120(x1120),
.x1121(x1121),
.x1122(x1122),
.x1123(x1123),
.x1124(x1124),
.x1125(x1125),
.x1126(x1126),
.x1127(x1127),
.x1128(x1128),
.x1129(x1129),
.x1130(x1130),
.x1131(x1131),
.x1132(x1132),
.x1133(x1133),
.x1134(x1134),
.x1135(x1135),
.x1136(x1136),
.x1137(x1137),
.x1138(x1138),
.x1139(x1139),
.x1140(x1140),
.x1141(x1141),
.x1142(x1142),
.x1143(x1143),
.x1144(x1144),
.x1145(x1145),
.x1146(x1146),
.x1147(x1147),
.x1148(x1148),
.x1149(x1149),
.x1150(x1150),
.x1151(x1151),
.x1152(x1152),
.x1153(x1153),
.x1154(x1154),
.x1155(x1155),
.x1156(x1156),
.x1157(x1157),
.x1158(x1158),
.x1159(x1159),
.x1160(x1160),
.x1161(x1161),
.x1162(x1162),
.x1163(x1163),
.x1164(x1164),
.x1165(x1165),
.x1166(x1166),
.x1167(x1167),
.x1168(x1168),
.x1169(x1169),
.x1170(x1170),
.x1171(x1171),
.x1172(x1172),
.x1173(x1173),
.x1174(x1174),
.x1175(x1175),
.x1176(x1176),
.x1177(x1177),
.x1178(x1178),
.x1179(x1179),
.x1180(x1180),
.x1181(x1181),
.x1182(x1182),
.x1183(x1183),
.x1184(x1184),
.x1185(x1185),
.x1186(x1186),
.x1187(x1187),
.x1188(x1188),
.x1189(x1189),
.x1190(x1190),
.x1191(x1191),
.x1192(x1192),
.x1193(x1193),
.x1194(x1194),
.x1195(x1195),
.x1196(x1196),
.x1197(x1197),
.x1198(x1198),
.x1199(x1199),
.x1200(x1200),
.x1201(x1201),
.x1202(x1202),
.x1203(x1203),
.x1204(x1204),
.x1205(x1205),
.x1206(x1206),
.x1207(x1207),
.x1208(x1208),
.x1209(x1209),
.x1210(x1210),
.x1211(x1211),
.x1212(x1212),
.x1213(x1213),
.x1214(x1214),
.x1215(x1215),
.x1216(x1216),
.x1217(x1217),
.x1218(x1218),
.x1219(x1219),
.x1220(x1220),
.x1221(x1221),
.x1222(x1222),
.x1223(x1223),
.x1224(x1224),
.x1225(x1225),
.x1226(x1226),
.x1227(x1227),
.x1228(x1228),
.x1229(x1229),
.x1230(x1230),
.x1231(x1231),
.x1232(x1232),
.x1233(x1233),
.x1234(x1234),
.x1235(x1235),
.x1236(x1236),
.x1237(x1237),
.x1238(x1238),
.x1239(x1239),
.x1240(x1240),
.x1241(x1241),
.x1242(x1242),
.x1243(x1243),
.x1244(x1244),
.x1245(x1245),
.x1246(x1246),
.x1247(x1247),
.x1248(x1248),
.x1249(x1249),
.x1250(x1250),
.x1251(x1251),
.x1252(x1252),
.x1253(x1253),
.x1254(x1254),
.x1255(x1255),
.x1256(x1256),
.x1257(x1257),
.x1258(x1258),
.x1259(x1259),
.x1260(x1260),
.x1261(x1261),
.x1262(x1262),
.x1263(x1263),
.x1264(x1264),
.x1265(x1265),
.x1266(x1266),
.x1267(x1267),
.x1268(x1268),
.x1269(x1269),
.x1270(x1270),
.x1271(x1271),
.x1272(x1272),
.x1273(x1273),
.x1274(x1274),
.x1275(x1275),
.x1276(x1276),
.x1277(x1277),
.x1278(x1278),
.x1279(x1279),
.x1280(x1280),
.x1281(x1281),
.x1282(x1282),
.x1283(x1283),
.x1284(x1284),
.x1285(x1285),
.x1286(x1286),
.x1287(x1287),
.x1288(x1288),
.x1289(x1289),
.x1290(x1290),
.x1291(x1291),
.x1292(x1292),
.x1293(x1293),
.x1294(x1294),
.x1295(x1295),
.x1296(x1296),
.x1297(x1297),
.x1298(x1298),
.x1299(x1299),
.x1300(x1300),
.x1301(x1301),
.x1302(x1302),
.x1303(x1303),
.x1304(x1304),
.x1305(x1305),
.x1306(x1306),
.x1307(x1307),
.x1308(x1308),
.x1309(x1309),
.x1310(x1310),
.x1311(x1311),
.x1312(x1312),
.x1313(x1313),
.x1314(x1314),
.x1315(x1315),
.x1316(x1316),
.x1317(x1317),
.x1318(x1318),
.x1319(x1319),
.x1320(x1320),
.x1321(x1321),
.x1322(x1322),
.x1323(x1323),
.x1324(x1324),
.x1325(x1325),
.x1326(x1326),
.x1327(x1327),
.x1328(x1328),
.x1329(x1329),
.x1330(x1330),
.x1331(x1331),
.x1332(x1332),
.x1333(x1333),
.x1334(x1334),
.x1335(x1335),
.x1336(x1336),
.x1337(x1337),
.x1338(x1338),
.x1339(x1339),
.x1340(x1340),
.x1341(x1341),
.x1342(x1342),
.x1343(x1343),
.x1344(x1344),
.x1345(x1345),
.x1346(x1346),
.x1347(x1347),
.x1348(x1348),
.x1349(x1349),
.x1350(x1350),
.x1351(x1351),
.x1352(x1352),
.x1353(x1353),
.x1354(x1354),
.x1355(x1355),
.x1356(x1356),
.x1357(x1357),
.x1358(x1358),
.x1359(x1359),
.x1360(x1360),
.x1361(x1361),
.x1362(x1362),
.x1363(x1363),
.x1364(x1364),
.x1365(x1365),
.x1366(x1366),
.x1367(x1367),
.x1368(x1368),
.x1369(x1369),
.x1370(x1370),
.x1371(x1371),
.x1372(x1372),
.x1373(x1373),
.x1374(x1374),
.x1375(x1375),
.x1376(x1376),
.x1377(x1377),
.x1378(x1378),
.x1379(x1379),
.x1380(x1380),
.x1381(x1381),
.x1382(x1382),
.x1383(x1383),
.x1384(x1384),
.x1385(x1385),
.x1386(x1386),
.x1387(x1387),
.x1388(x1388),
.x1389(x1389),
.x1390(x1390),
.x1391(x1391),
.x1392(x1392),
.x1393(x1393),
.x1394(x1394),
.x1395(x1395),
.x1396(x1396),
.x1397(x1397),
.x1398(x1398),
.x1399(x1399),
.x1400(x1400),
.x1401(x1401),
.x1402(x1402),
.x1403(x1403),
.x1404(x1404),
.x1405(x1405),
.x1406(x1406),
.x1407(x1407),
.x1408(x1408),
.x1409(x1409),
.x1410(x1410),
.x1411(x1411),
.x1412(x1412),
.x1413(x1413),
.x1414(x1414),
.x1415(x1415),
.x1416(x1416),
.x1417(x1417),
.x1418(x1418),
.x1419(x1419),
.x1420(x1420),
.x1421(x1421),
.x1422(x1422),
.x1423(x1423),
.x1424(x1424),
.x1425(x1425),
.x1426(x1426),
.x1427(x1427),
.x1428(x1428),
.x1429(x1429),
.x1430(x1430),
.x1431(x1431),
.x1432(x1432),
.x1433(x1433),
.x1434(x1434),
.x1435(x1435),
.x1436(x1436),
.x1437(x1437),
.x1438(x1438),
.x1439(x1439),
.x1440(x1440),
.x1441(x1441),
.x1442(x1442),
.x1443(x1443),
.x1444(x1444),
.x1445(x1445),
.x1446(x1446),
.x1447(x1447),
.x1448(x1448),
.x1449(x1449),
.x1450(x1450),
.x1451(x1451),
.x1452(x1452),
.x1453(x1453),
.x1454(x1454),
.x1455(x1455),
.x1456(x1456),
.x1457(x1457),
.x1458(x1458),
.x1459(x1459),
.x1460(x1460),
.x1461(x1461),
.x1462(x1462),
.x1463(x1463),
.x1464(x1464),
.x1465(x1465),
.x1466(x1466),
.x1467(x1467),
.x1468(x1468),
.x1469(x1469),
.x1470(x1470),
.x1471(x1471),
.x1472(x1472),
.x1473(x1473),
.x1474(x1474),
.x1475(x1475),
.x1476(x1476),
.x1477(x1477),
.x1478(x1478),
.x1479(x1479),
.x1480(x1480),
.x1481(x1481),
.x1482(x1482),
.x1483(x1483),
.x1484(x1484),
.x1485(x1485),
.x1486(x1486),
.x1487(x1487),
.x1488(x1488),
.x1489(x1489),
.x1490(x1490),
.x1491(x1491),
.x1492(x1492),
.x1493(x1493),
.x1494(x1494),
.x1495(x1495),
.x1496(x1496),
.x1497(x1497),
.x1498(x1498),
.x1499(x1499),
.x1500(x1500),
.x1501(x1501),
.x1502(x1502),
.x1503(x1503),
.x1504(x1504),
.x1505(x1505),
.x1506(x1506),
.x1507(x1507),
.x1508(x1508),
.x1509(x1509),
.x1510(x1510),
.x1511(x1511),
.x1512(x1512),
.x1513(x1513),
.x1514(x1514),
.x1515(x1515),
.x1516(x1516),
.x1517(x1517),
.x1518(x1518),
.x1519(x1519),
.x1520(x1520),
.x1521(x1521),
.x1522(x1522),
.x1523(x1523),
.x1524(x1524),
.x1525(x1525),
.x1526(x1526),
.x1527(x1527),
.x1528(x1528),
.x1529(x1529),
.x1530(x1530),
.x1531(x1531),
.x1532(x1532),
.x1533(x1533),
.x1534(x1534),
.x1535(x1535),
.x1536(x1536),
.x1537(x1537),
.x1538(x1538),
.x1539(x1539),
.x1540(x1540),
.x1541(x1541),
.x1542(x1542),
.x1543(x1543),
.x1544(x1544),
.x1545(x1545),
.x1546(x1546),
.x1547(x1547),
.x1548(x1548),
.x1549(x1549),
.x1550(x1550),
.x1551(x1551),
.x1552(x1552),
.x1553(x1553),
.x1554(x1554),
.x1555(x1555),
.x1556(x1556),
.x1557(x1557),
.x1558(x1558),
.x1559(x1559),
.x1560(x1560),
.x1561(x1561),
.x1562(x1562),
.x1563(x1563),
.x1564(x1564),
.x1565(x1565),
.x1566(x1566),
.x1567(x1567),
.x1568(x1568),
.x1569(x1569),
.x1570(x1570),
.x1571(x1571),
.x1572(x1572),
.x1573(x1573),
.x1574(x1574),
.x1575(x1575),
.x1576(x1576),
.x1577(x1577),
.x1578(x1578),
.x1579(x1579),
.x1580(x1580),
.x1581(x1581),
.x1582(x1582),
.x1583(x1583),
.x1584(x1584),
.x1585(x1585),
.x1586(x1586),
.x1587(x1587),
.x1588(x1588),
.x1589(x1589),
.x1590(x1590),
.x1591(x1591),
.x1592(x1592),
.x1593(x1593),
.x1594(x1594),
.x1595(x1595),
.x1596(x1596),
.x1597(x1597),
.x1598(x1598),
.x1599(x1599),
.x1600(x1600),
.x1601(x1601),
.x1602(x1602),
.x1603(x1603),
.x1604(x1604),
.x1605(x1605),
.x1606(x1606),
.x1607(x1607),
.x1608(x1608),
.x1609(x1609),
.x1610(x1610),
.x1611(x1611),
.x1612(x1612),
.x1613(x1613),
.x1614(x1614),
.x1615(x1615),
.x1616(x1616),
.x1617(x1617),
.x1618(x1618),
.x1619(x1619),
.x1620(x1620),
.x1621(x1621),
.x1622(x1622),
.x1623(x1623),
.x1624(x1624),
.x1625(x1625),
.x1626(x1626),
.x1627(x1627),
.x1628(x1628),
.x1629(x1629),
.x1630(x1630),
.x1631(x1631),
.x1632(x1632),
.x1633(x1633),
.x1634(x1634),
.x1635(x1635),
.x1636(x1636),
.x1637(x1637),
.x1638(x1638),
.x1639(x1639),
.x1640(x1640),
.x1641(x1641),
.x1642(x1642),
.x1643(x1643),
.x1644(x1644),
.x1645(x1645),
.x1646(x1646),
.x1647(x1647),
.x1648(x1648),
.x1649(x1649),
.x1650(x1650),
.x1651(x1651),
.x1652(x1652),
.x1653(x1653),
.x1654(x1654),
.x1655(x1655),
.x1656(x1656),
.x1657(x1657),
.x1658(x1658),
.x1659(x1659),
.x1660(x1660),
.x1661(x1661),
.x1662(x1662),
.x1663(x1663),
.x1664(x1664),
.x1665(x1665),
.x1666(x1666),
.x1667(x1667),
.x1668(x1668),
.x1669(x1669),
.x1670(x1670),
.x1671(x1671),
.x1672(x1672),
.x1673(x1673),
.x1674(x1674),
.x1675(x1675),
.x1676(x1676),
.x1677(x1677),
.x1678(x1678),
.x1679(x1679),
.x1680(x1680),
.x1681(x1681),
.x1682(x1682),
.x1683(x1683),
.x1684(x1684),
.x1685(x1685),
.x1686(x1686),
.x1687(x1687),
.x1688(x1688),
.x1689(x1689),
.x1690(x1690),
.x1691(x1691),
.x1692(x1692),
.x1693(x1693),
.x1694(x1694),
.x1695(x1695),
.x1696(x1696),
.x1697(x1697),
.x1698(x1698),
.x1699(x1699),
.x1700(x1700),
.x1701(x1701),
.x1702(x1702),
.x1703(x1703),
.x1704(x1704),
.x1705(x1705),
.x1706(x1706),
.x1707(x1707),
.x1708(x1708),
.x1709(x1709),
.x1710(x1710),
.x1711(x1711),
.x1712(x1712),
.x1713(x1713),
.x1714(x1714),
.x1715(x1715),
.x1716(x1716),
.x1717(x1717),
.x1718(x1718),
.x1719(x1719),
.x1720(x1720),
.x1721(x1721),
.x1722(x1722),
.x1723(x1723),
.x1724(x1724),
.x1725(x1725),
.x1726(x1726),
.x1727(x1727),
.x1728(x1728),
.x1729(x1729),
.x1730(x1730),
.x1731(x1731),
.x1732(x1732),
.x1733(x1733),
.x1734(x1734),
.x1735(x1735),
.x1736(x1736),
.x1737(x1737),
.x1738(x1738),
.x1739(x1739),
.x1740(x1740),
.x1741(x1741),
.x1742(x1742),
.x1743(x1743),
.x1744(x1744),
.x1745(x1745),
.x1746(x1746),
.x1747(x1747),
.x1748(x1748),
.x1749(x1749),
.x1750(x1750),
.x1751(x1751),
.x1752(x1752),
.x1753(x1753),
.x1754(x1754),
.x1755(x1755),
.x1756(x1756),
.x1757(x1757),
.x1758(x1758),
.x1759(x1759),
.x1760(x1760),
.x1761(x1761),
.x1762(x1762),
.x1763(x1763),
.x1764(x1764),
.x1765(x1765),
.x1766(x1766),
.x1767(x1767),
.x1768(x1768),
.x1769(x1769),
.x1770(x1770),
.x1771(x1771),
.x1772(x1772),
.x1773(x1773),
.x1774(x1774),
.x1775(x1775),
.x1776(x1776),
.x1777(x1777),
.x1778(x1778),
.x1779(x1779),
.x1780(x1780),
.x1781(x1781),
.x1782(x1782),
.x1783(x1783),
.x1784(x1784),
.x1785(x1785),
.x1786(x1786),
.x1787(x1787),
.x1788(x1788),
.x1789(x1789),
.x1790(x1790),
.x1791(x1791),
.x1792(x1792),
.x1793(x1793),
.x1794(x1794),
.x1795(x1795),
.x1796(x1796),
.x1797(x1797),
.x1798(x1798),
.x1799(x1799),
.x1800(x1800),
.x1801(x1801),
.x1802(x1802),
.x1803(x1803),
.x1804(x1804),
.x1805(x1805),
.x1806(x1806),
.x1807(x1807),
.x1808(x1808),
.x1809(x1809),
.x1810(x1810),
.x1811(x1811),
.x1812(x1812),
.x1813(x1813),
.x1814(x1814),
.x1815(x1815),
.x1816(x1816),
.x1817(x1817),
.x1818(x1818),
.x1819(x1819),
.x1820(x1820),
.x1821(x1821),
.x1822(x1822),
.x1823(x1823),
.x1824(x1824),
.x1825(x1825),
.x1826(x1826),
.x1827(x1827),
.x1828(x1828),
.x1829(x1829),
.x1830(x1830),
.x1831(x1831),
.x1832(x1832),
.x1833(x1833),
.x1834(x1834),
.x1835(x1835),
.x1836(x1836),
.x1837(x1837),
.x1838(x1838),
.x1839(x1839),
.x1840(x1840),
.x1841(x1841),
.x1842(x1842),
.x1843(x1843),
.x1844(x1844),
.x1845(x1845),
.x1846(x1846),
.x1847(x1847),
.x1848(x1848),
.x1849(x1849),
.x1850(x1850),
.x1851(x1851),
.x1852(x1852),
.x1853(x1853),
.x1854(x1854),
.x1855(x1855),
.x1856(x1856),
.x1857(x1857),
.x1858(x1858),
.x1859(x1859),
.x1860(x1860),
.x1861(x1861),
.x1862(x1862),
.x1863(x1863),
.x1864(x1864),
.x1865(x1865),
.x1866(x1866),
.x1867(x1867),
.x1868(x1868),
.x1869(x1869),
.x1870(x1870),
.x1871(x1871),
.x1872(x1872),
.x1873(x1873),
.x1874(x1874),
.x1875(x1875),
.x1876(x1876),
.x1877(x1877),
.x1878(x1878),
.x1879(x1879),
.x1880(x1880),
.x1881(x1881),
.x1882(x1882),
.x1883(x1883),
.x1884(x1884),
.x1885(x1885),
.x1886(x1886),
.x1887(x1887),
.x1888(x1888),
.x1889(x1889),
.x1890(x1890),
.x1891(x1891),
.x1892(x1892),
.x1893(x1893),
.x1894(x1894),
.x1895(x1895),
.x1896(x1896),
.x1897(x1897),
.x1898(x1898),
.x1899(x1899),
.x1900(x1900),
.x1901(x1901),
.x1902(x1902),
.x1903(x1903),
.x1904(x1904),
.x1905(x1905),
.x1906(x1906),
.x1907(x1907),
.x1908(x1908),
.x1909(x1909),
.x1910(x1910),
.x1911(x1911),
.x1912(x1912),
.x1913(x1913),
.x1914(x1914),
.x1915(x1915),
.x1916(x1916),
.x1917(x1917),
.x1918(x1918),
.x1919(x1919),
.x1920(x1920),
.x1921(x1921),
.x1922(x1922),
.x1923(x1923),
.x1924(x1924),
.x1925(x1925),
.x1926(x1926),
.x1927(x1927),
.x1928(x1928),
.x1929(x1929),
.x1930(x1930),
.x1931(x1931),
.x1932(x1932),
.x1933(x1933),
.x1934(x1934),
.x1935(x1935),
.x1936(x1936),
.x1937(x1937),
.x1938(x1938),
.x1939(x1939),
.x1940(x1940),
.x1941(x1941),
.x1942(x1942),
.x1943(x1943),
.x1944(x1944),
.x1945(x1945),
.x1946(x1946),
.x1947(x1947),
.x1948(x1948),
.x1949(x1949),
.x1950(x1950),
.x1951(x1951),
.x1952(x1952),
.x1953(x1953),
.x1954(x1954),
.x1955(x1955),
.x1956(x1956),
.x1957(x1957),
.x1958(x1958),
.x1959(x1959),
.x1960(x1960),
.x1961(x1961),
.x1962(x1962),
.x1963(x1963),
.x1964(x1964),
.x1965(x1965),
.x1966(x1966),
.x1967(x1967),
.x1968(x1968),
.x1969(x1969),
.x1970(x1970),
.x1971(x1971),
.x1972(x1972),
.x1973(x1973),
.x1974(x1974),
.x1975(x1975),
.x1976(x1976),
.x1977(x1977),
.x1978(x1978),
.x1979(x1979),
.x1980(x1980),
.x1981(x1981),
.x1982(x1982),
.x1983(x1983),
.x1984(x1984),
.x1985(x1985),
.x1986(x1986),
.x1987(x1987),
.x1988(x1988),
.x1989(x1989),
.x1990(x1990),
.x1991(x1991),
.x1992(x1992),
.x1993(x1993),
.x1994(x1994),
.x1995(x1995),
.x1996(x1996),
.x1997(x1997),
.x1998(x1998),
.x1999(x1999),
.x2000(x2000),
.x2001(x2001),
.x2002(x2002),
.x2003(x2003),
.x2004(x2004),
.x2005(x2005),
.x2006(x2006),
.x2007(x2007),
.x2008(x2008),
.x2009(x2009),
.x2010(x2010),
.x2011(x2011),
.x2012(x2012),
.x2013(x2013),
.x2014(x2014),
.x2015(x2015),
.x2016(x2016),
.x2017(x2017),
.x2018(x2018),
.x2019(x2019),
.x2020(x2020),
.x2021(x2021),
.x2022(x2022),
.x2023(x2023),
.x2024(x2024),
.x2025(x2025),
.x2026(x2026),
.x2027(x2027),
.x2028(x2028),
.x2029(x2029),
.x2030(x2030),
.x2031(x2031),
.x2032(x2032),
.x2033(x2033),
.x2034(x2034),
.x2035(x2035),
.x2036(x2036),
.x2037(x2037),
.x2038(x2038),
.x2039(x2039),
.x2040(x2040),
.x2041(x2041),
.x2042(x2042),
.x2043(x2043),
.x2044(x2044),
.x2045(x2045),
.x2046(x2046),
.x2047(x2047),
.x2048(x2048),
.x2049(x2049),
.x2050(x2050),
.x2051(x2051),
.x2052(x2052),
.x2053(x2053),
.x2054(x2054),
.x2055(x2055),
.x2056(x2056),
.x2057(x2057),
.x2058(x2058),
.x2059(x2059),
.x2060(x2060),
.x2061(x2061),
.x2062(x2062),
.x2063(x2063),
.x2064(x2064),
.x2065(x2065),
.x2066(x2066),
.x2067(x2067),
.x2068(x2068),
.x2069(x2069),
.x2070(x2070),
.x2071(x2071),
.x2072(x2072),
.x2073(x2073),
.x2074(x2074),
.x2075(x2075),
.x2076(x2076),
.x2077(x2077),
.x2078(x2078),
.x2079(x2079),
.x2080(x2080),
.x2081(x2081),
.x2082(x2082),
.x2083(x2083),
.x2084(x2084),
.x2085(x2085),
.x2086(x2086),
.x2087(x2087),
.x2088(x2088),
.x2089(x2089),
.x2090(x2090),
.x2091(x2091),
.x2092(x2092),
.x2093(x2093),
.x2094(x2094),
.x2095(x2095),
.x2096(x2096),
.x2097(x2097),
.x2098(x2098),
.x2099(x2099),
.x2100(x2100),
.x2101(x2101),
.x2102(x2102),
.x2103(x2103),
.x2104(x2104),
.x2105(x2105),
.x2106(x2106),
.x2107(x2107),
.x2108(x2108),
.x2109(x2109),
.x2110(x2110),
.x2111(x2111),
.x2112(x2112),
.x2113(x2113),
.x2114(x2114),
.x2115(x2115),
.x2116(x2116),
.x2117(x2117),
.x2118(x2118),
.x2119(x2119),
.x2120(x2120),
.x2121(x2121),
.x2122(x2122),
.x2123(x2123),
.x2124(x2124),
.x2125(x2125),
.x2126(x2126),
.x2127(x2127),
.x2128(x2128),
.x2129(x2129),
.x2130(x2130),
.x2131(x2131),
.x2132(x2132),
.x2133(x2133),
.x2134(x2134),
.x2135(x2135),
.x2136(x2136),
.x2137(x2137),
.x2138(x2138),
.x2139(x2139),
.x2140(x2140),
.x2141(x2141),
.x2142(x2142),
.x2143(x2143),
.x2144(x2144),
.x2145(x2145),
.x2146(x2146),
.x2147(x2147),
.x2148(x2148),
.x2149(x2149),
.x2150(x2150),
.x2151(x2151),
.x2152(x2152),
.x2153(x2153),
.x2154(x2154),
.x2155(x2155),
.x2156(x2156),
.x2157(x2157),
.x2158(x2158),
.x2159(x2159),
.x2160(x2160),
.x2161(x2161),
.x2162(x2162),
.x2163(x2163),
.x2164(x2164),
.x2165(x2165),
.x2166(x2166),
.x2167(x2167),
.x2168(x2168),
.x2169(x2169),
.x2170(x2170),
.x2171(x2171),
.x2172(x2172),
.x2173(x2173),
.x2174(x2174),
.x2175(x2175),
.x2176(x2176),
.x2177(x2177),
.x2178(x2178),
.x2179(x2179),
.x2180(x2180),
.x2181(x2181),
.x2182(x2182),
.x2183(x2183),
.x2184(x2184),
.x2185(x2185),
.x2186(x2186),
.x2187(x2187),
.x2188(x2188),
.x2189(x2189),
.x2190(x2190),
.x2191(x2191),
.x2192(x2192),
.x2193(x2193),
.x2194(x2194),
.x2195(x2195),
.x2196(x2196),
.x2197(x2197),
.x2198(x2198),
.x2199(x2199),
.x2200(x2200),
.x2201(x2201),
.x2202(x2202),
.x2203(x2203),
.x2204(x2204),
.x2205(x2205),
.x2206(x2206),
.x2207(x2207),
.x2208(x2208),
.x2209(x2209),
.x2210(x2210),
.x2211(x2211),
.x2212(x2212),
.x2213(x2213),
.x2214(x2214),
.x2215(x2215),
.x2216(x2216),
.x2217(x2217),
.x2218(x2218),
.x2219(x2219),
.x2220(x2220),
.x2221(x2221),
.x2222(x2222),
.x2223(x2223),
.x2224(x2224),
.x2225(x2225),
.x2226(x2226),
.x2227(x2227),
.x2228(x2228),
.x2229(x2229),
.x2230(x2230),
.x2231(x2231),
.x2232(x2232),
.x2233(x2233),
.x2234(x2234),
.x2235(x2235),
.x2236(x2236),
.x2237(x2237),
.x2238(x2238),
.x2239(x2239),
.x2240(x2240),
.x2241(x2241),
.x2242(x2242),
.x2243(x2243),
.x2244(x2244),
.x2245(x2245),
.x2246(x2246),
.x2247(x2247),
.x2248(x2248),
.x2249(x2249),
.x2250(x2250),
.x2251(x2251),
.x2252(x2252),
.x2253(x2253),
.x2254(x2254),
.x2255(x2255),
.x2256(x2256),
.x2257(x2257),
.x2258(x2258),
.x2259(x2259),
.x2260(x2260),
.x2261(x2261),
.x2262(x2262),
.x2263(x2263),
.x2264(x2264),
.x2265(x2265),
.x2266(x2266),
.x2267(x2267),
.x2268(x2268),
.x2269(x2269),
.x2270(x2270),
.x2271(x2271),
.x2272(x2272),
.x2273(x2273),
.x2274(x2274),
.x2275(x2275),
.x2276(x2276),
.x2277(x2277),
.x2278(x2278),
.x2279(x2279),
.x2280(x2280),
.x2281(x2281),
.x2282(x2282),
.x2283(x2283),
.x2284(x2284),
.x2285(x2285),
.x2286(x2286),
.x2287(x2287),
.x2288(x2288),
.x2289(x2289),
.x2290(x2290),
.x2291(x2291),
.x2292(x2292),
.x2293(x2293),
.x2294(x2294),
.x2295(x2295),
.x2296(x2296),
.x2297(x2297),
.x2298(x2298),
.x2299(x2299),
.x2300(x2300),
.x2301(x2301),
.x2302(x2302),
.x2303(x2303),
.x2304(x2304),
.x2305(x2305),
.x2306(x2306),
.x2307(x2307),
.x2308(x2308),
.x2309(x2309),
.x2310(x2310),
.x2311(x2311),
.x2312(x2312),
.x2313(x2313),
.x2314(x2314),
.x2315(x2315),
.x2316(x2316),
.x2317(x2317),
.x2318(x2318),
.x2319(x2319),
.x2320(x2320),
.x2321(x2321),
.x2322(x2322),
.x2323(x2323),
.x2324(x2324),
.x2325(x2325),
.x2326(x2326),
.x2327(x2327),
.x2328(x2328),
.x2329(x2329),
.x2330(x2330),
.x2331(x2331),
.x2332(x2332),
.x2333(x2333),
.x2334(x2334),
.x2335(x2335),
.x2336(x2336),
.x2337(x2337),
.x2338(x2338),
.x2339(x2339),
.x2340(x2340),
.x2341(x2341),
.x2342(x2342),
.x2343(x2343),
.x2344(x2344),
.x2345(x2345),
.x2346(x2346),
.x2347(x2347),
.x2348(x2348),
.x2349(x2349),
.x2350(x2350),
.x2351(x2351),
.x2352(x2352),
.x2353(x2353),
.x2354(x2354),
.x2355(x2355),
.x2356(x2356),
.x2357(x2357),
.x2358(x2358),
.x2359(x2359),
.x2360(x2360),
.x2361(x2361),
.x2362(x2362),
.x2363(x2363),
.x2364(x2364),
.x2365(x2365),
.x2366(x2366),
.x2367(x2367),
.x2368(x2368),
.x2369(x2369),
.x2370(x2370),
.x2371(x2371),
.x2372(x2372),
.x2373(x2373),
.x2374(x2374),
.x2375(x2375),
.x2376(x2376),
.x2377(x2377),
.x2378(x2378),
.x2379(x2379),
.x2380(x2380),
.x2381(x2381),
.x2382(x2382),
.x2383(x2383),
.x2384(x2384),
.x2385(x2385),
.x2386(x2386),
.x2387(x2387),
.x2388(x2388),
.x2389(x2389),
.x2390(x2390),
.x2391(x2391),
.x2392(x2392),
.x2393(x2393),
.x2394(x2394),
.x2395(x2395),
.x2396(x2396),
.x2397(x2397),
.x2398(x2398),
.x2399(x2399),
.x2400(x2400),
.x2401(x2401),
.x2402(x2402),
.x2403(x2403),
.x2404(x2404),
.x2405(x2405),
.x2406(x2406),
.x2407(x2407),
.x2408(x2408),
.x2409(x2409),
.x2410(x2410),
.x2411(x2411),
.x2412(x2412),
.x2413(x2413),
.x2414(x2414),
.x2415(x2415),
.x2416(x2416),
.x2417(x2417),
.x2418(x2418),
.x2419(x2419),
.x2420(x2420),
.x2421(x2421),
.x2422(x2422),
.x2423(x2423),
.x2424(x2424),
.x2425(x2425),
.x2426(x2426),
.x2427(x2427),
.x2428(x2428),
.x2429(x2429),
.x2430(x2430),
.x2431(x2431),
.x2432(x2432),
.x2433(x2433),
.x2434(x2434),
.x2435(x2435),
.x2436(x2436),
.x2437(x2437),
.x2438(x2438),
.x2439(x2439),
.x2440(x2440),
.x2441(x2441),
.x2442(x2442),
.x2443(x2443),
.x2444(x2444),
.x2445(x2445),
.x2446(x2446),
.x2447(x2447),
.x2448(x2448),
.x2449(x2449),
.x2450(x2450),
.x2451(x2451),
.x2452(x2452),
.x2453(x2453),
.x2454(x2454),
.x2455(x2455),
.x2456(x2456),
.x2457(x2457),
.x2458(x2458),
.x2459(x2459),
.x2460(x2460),
.x2461(x2461),
.x2462(x2462),
.x2463(x2463),
.x2464(x2464),
.x2465(x2465),
.x2466(x2466),
.x2467(x2467),
.x2468(x2468),
.x2469(x2469),
.x2470(x2470),
.x2471(x2471),
.x2472(x2472),
.x2473(x2473),
.x2474(x2474),
.x2475(x2475),
.x2476(x2476),
.x2477(x2477),
.x2478(x2478),
.x2479(x2479),
.x2480(x2480),
.x2481(x2481),
.x2482(x2482),
.x2483(x2483),
.x2484(x2484),
.x2485(x2485),
.x2486(x2486),
.x2487(x2487),
.x2488(x2488),
.x2489(x2489),
.x2490(x2490),
.x2491(x2491),
.x2492(x2492),
.x2493(x2493),
.x2494(x2494),
.x2495(x2495),
.x2496(x2496),
.x2497(x2497),
.x2498(x2498),
.x2499(x2499),
.x2500(x2500),
.x2501(x2501),
.x2502(x2502),
.x2503(x2503),
.x2504(x2504),
.x2505(x2505),
.x2506(x2506),
.x2507(x2507),
.x2508(x2508),
.x2509(x2509),
.x2510(x2510),
.x2511(x2511),
.x2512(x2512),
.x2513(x2513),
.x2514(x2514),
.x2515(x2515),
.x2516(x2516),
.x2517(x2517),
.x2518(x2518),
.x2519(x2519),
.x2520(x2520),
.x2521(x2521),
.x2522(x2522),
.x2523(x2523),
.x2524(x2524),
.x2525(x2525),
.x2526(x2526),
.x2527(x2527),
.x2528(x2528),
.x2529(x2529),
.x2530(x2530),
.x2531(x2531),
.x2532(x2532),
.x2533(x2533),
.x2534(x2534),
.x2535(x2535),
.x2536(x2536),
.x2537(x2537),
.x2538(x2538),
.x2539(x2539),
.x2540(x2540),
.x2541(x2541),
.x2542(x2542),
.x2543(x2543),
.x2544(x2544),
.x2545(x2545),
.x2546(x2546),
.x2547(x2547),
.x2548(x2548),
.x2549(x2549),
.x2550(x2550),
.x2551(x2551),
.x2552(x2552),
.x2553(x2553),
.x2554(x2554),
.x2555(x2555),
.x2556(x2556),
.x2557(x2557),
.x2558(x2558),
.x2559(x2559),
.x2560(x2560),
.x2561(x2561),
.x2562(x2562),
.x2563(x2563),
.x2564(x2564),
.x2565(x2565),
.x2566(x2566),
.x2567(x2567),
.x2568(x2568),
.x2569(x2569),
.x2570(x2570),
.x2571(x2571),
.x2572(x2572),
.x2573(x2573),
.x2574(x2574),
.x2575(x2575),
.x2576(x2576),
.x2577(x2577),
.x2578(x2578),
.x2579(x2579),
.x2580(x2580),
.x2581(x2581),
.x2582(x2582),
.x2583(x2583),
.x2584(x2584),
.x2585(x2585),
.x2586(x2586),
.x2587(x2587),
.x2588(x2588),
.x2589(x2589),
.x2590(x2590),
.x2591(x2591),
.x2592(x2592),
.x2593(x2593),
.x2594(x2594),
.x2595(x2595),
.x2596(x2596),
.x2597(x2597),
.x2598(x2598),
.x2599(x2599),
.x2600(x2600),
.x2601(x2601),
.x2602(x2602),
.x2603(x2603),
.x2604(x2604),
.x2605(x2605),
.x2606(x2606),
.x2607(x2607),
.x2608(x2608),
.x2609(x2609),
.x2610(x2610),
.x2611(x2611),
.x2612(x2612),
.x2613(x2613),
.x2614(x2614),
.x2615(x2615),
.x2616(x2616),
.x2617(x2617),
.x2618(x2618),
.x2619(x2619),
.x2620(x2620),
.x2621(x2621),
.x2622(x2622),
.x2623(x2623),
.x2624(x2624),
.x2625(x2625),
.x2626(x2626),
.x2627(x2627),
.x2628(x2628),
.x2629(x2629),
.x2630(x2630),
.x2631(x2631),
.x2632(x2632),
.x2633(x2633),
.x2634(x2634),
.x2635(x2635),
.x2636(x2636),
.x2637(x2637),
.x2638(x2638),
.x2639(x2639),
.x2640(x2640),
.x2641(x2641),
.x2642(x2642),
.x2643(x2643),
.x2644(x2644),
.x2645(x2645),
.x2646(x2646),
.x2647(x2647),
.x2648(x2648),
.x2649(x2649),
.x2650(x2650),
.x2651(x2651),
.x2652(x2652),
.x2653(x2653),
.x2654(x2654),
.x2655(x2655),
.x2656(x2656),
.x2657(x2657),
.x2658(x2658),
.x2659(x2659),
.x2660(x2660),
.x2661(x2661),
.x2662(x2662),
.x2663(x2663),
.x2664(x2664),
.x2665(x2665),
.x2666(x2666),
.x2667(x2667),
.x2668(x2668),
.x2669(x2669),
.x2670(x2670),
.x2671(x2671),
.x2672(x2672),
.x2673(x2673),
.x2674(x2674),
.x2675(x2675),
.x2676(x2676),
.x2677(x2677),
.x2678(x2678),
.x2679(x2679),
.x2680(x2680),
.x2681(x2681),
.x2682(x2682),
.x2683(x2683),
.x2684(x2684),
.x2685(x2685),
.x2686(x2686),
.x2687(x2687),
.x2688(x2688),
.x2689(x2689),
.x2690(x2690),
.x2691(x2691),
.x2692(x2692),
.x2693(x2693),
.x2694(x2694),
.x2695(x2695),
.x2696(x2696),
.x2697(x2697),
.x2698(x2698),
.x2699(x2699),
.x2700(x2700),
.x2701(x2701),
.x2702(x2702),
.x2703(x2703),
.x2704(x2704),
.x2705(x2705),
.x2706(x2706),
.x2707(x2707),
.x2708(x2708),
.x2709(x2709),
.x2710(x2710),
.x2711(x2711),
.x2712(x2712),
.x2713(x2713),
.x2714(x2714),
.x2715(x2715),
.x2716(x2716),
.x2717(x2717),
.x2718(x2718),
.x2719(x2719),
.x2720(x2720),
.x2721(x2721),
.x2722(x2722),
.x2723(x2723),
.x2724(x2724),
.x2725(x2725),
.x2726(x2726),
.x2727(x2727),
.x2728(x2728),
.x2729(x2729),
.x2730(x2730),
.x2731(x2731),
.x2732(x2732),
.x2733(x2733),
.x2734(x2734),
.x2735(x2735),
.x2736(x2736),
.x2737(x2737),
.x2738(x2738),
.x2739(x2739),
.x2740(x2740),
.x2741(x2741),
.x2742(x2742),
.x2743(x2743),
.x2744(x2744),
.x2745(x2745),
.x2746(x2746),
.x2747(x2747),
.x2748(x2748),
.x2749(x2749),
.x2750(x2750),
.x2751(x2751),
.x2752(x2752),
.x2753(x2753),
.x2754(x2754),
.x2755(x2755),
.x2756(x2756),
.x2757(x2757),
.x2758(x2758),
.x2759(x2759),
.x2760(x2760),
.x2761(x2761),
.x2762(x2762),
.x2763(x2763),
.x2764(x2764),
.x2765(x2765),
.x2766(x2766),
.x2767(x2767),
.x2768(x2768),
.x2769(x2769),
.x2770(x2770),
.x2771(x2771),
.x2772(x2772),
.x2773(x2773),
.x2774(x2774),
.x2775(x2775),
.x2776(x2776),
.x2777(x2777),
.x2778(x2778),
.x2779(x2779),
.x2780(x2780),
.x2781(x2781),
.x2782(x2782),
.x2783(x2783),
.x2784(x2784),
.x2785(x2785),
.x2786(x2786),
.x2787(x2787),
.x2788(x2788),
.x2789(x2789),
.x2790(x2790),
.x2791(x2791),
.x2792(x2792),
.x2793(x2793),
.x2794(x2794),
.x2795(x2795),
.x2796(x2796),
.x2797(x2797),
.x2798(x2798),
.x2799(x2799),
.x2800(x2800),
.x2801(x2801),
.x2802(x2802),
.x2803(x2803),
.x2804(x2804),
.x2805(x2805),
.x2806(x2806),
.x2807(x2807),
.x2808(x2808),
.x2809(x2809),
.x2810(x2810),
.x2811(x2811),
.x2812(x2812),
.x2813(x2813),
.x2814(x2814),
.x2815(x2815),
.x2816(x2816),
.x2817(x2817),
.x2818(x2818),
.x2819(x2819),
.x2820(x2820),
.x2821(x2821),
.x2822(x2822),
.x2823(x2823),
.x2824(x2824),
.x2825(x2825),
.x2826(x2826),
.x2827(x2827),
.x2828(x2828),
.x2829(x2829),
.x2830(x2830),
.x2831(x2831),
.x2832(x2832),
.x2833(x2833),
.x2834(x2834),
.x2835(x2835),
.x2836(x2836),
.x2837(x2837),
.x2838(x2838),
.x2839(x2839),
.x2840(x2840),
.x2841(x2841),
.x2842(x2842),
.x2843(x2843),
.x2844(x2844),
.x2845(x2845),
.x2846(x2846),
.x2847(x2847),
.x2848(x2848),
.x2849(x2849),
.x2850(x2850),
.x2851(x2851),
.x2852(x2852),
.x2853(x2853),
.x2854(x2854),
.x2855(x2855),
.x2856(x2856),
.x2857(x2857),
.x2858(x2858),
.x2859(x2859),
.x2860(x2860),
.x2861(x2861),
.x2862(x2862),
.x2863(x2863),
.x2864(x2864),
.x2865(x2865),
.x2866(x2866),
.x2867(x2867),
.x2868(x2868),
.x2869(x2869),
.x2870(x2870),
.x2871(x2871),
.x2872(x2872),
.x2873(x2873),
.x2874(x2874),
.x2875(x2875),
.x2876(x2876),
.x2877(x2877),
.x2878(x2878),
.x2879(x2879),
.x2880(x2880),
.x2881(x2881),
.x2882(x2882),
.x2883(x2883),
.x2884(x2884),
.x2885(x2885),
.x2886(x2886),
.x2887(x2887),
.x2888(x2888),
.x2889(x2889),
.x2890(x2890),
.x2891(x2891),
.x2892(x2892),
.x2893(x2893),
.x2894(x2894),
.x2895(x2895),
.x2896(x2896),
.x2897(x2897),
.x2898(x2898),
.x2899(x2899),
.x2900(x2900),
.x2901(x2901),
.x2902(x2902),
.x2903(x2903),
.x2904(x2904),
.x2905(x2905),
.x2906(x2906),
.x2907(x2907),
.x2908(x2908),
.x2909(x2909),
.x2910(x2910),
.x2911(x2911),
.x2912(x2912),
.x2913(x2913),
.x2914(x2914),
.x2915(x2915),
.x2916(x2916),
.x2917(x2917),
.x2918(x2918),
.x2919(x2919),
.x2920(x2920),
.x2921(x2921),
.x2922(x2922),
.x2923(x2923),
.x2924(x2924),
.x2925(x2925),
.x2926(x2926),
.x2927(x2927),
.x2928(x2928),
.x2929(x2929),
.x2930(x2930),
.x2931(x2931),
.x2932(x2932),
.x2933(x2933),
.x2934(x2934),
.x2935(x2935),
.x2936(x2936),
.x2937(x2937),
.x2938(x2938),
.x2939(x2939),
.x2940(x2940),
.x2941(x2941),
.x2942(x2942),
.x2943(x2943),
.x2944(x2944),
.x2945(x2945),
.x2946(x2946),
.x2947(x2947),
.x2948(x2948),
.x2949(x2949),
.x2950(x2950),
.x2951(x2951),
.x2952(x2952),
.x2953(x2953),
.x2954(x2954),
.x2955(x2955),
.x2956(x2956),
.x2957(x2957),
.x2958(x2958),
.x2959(x2959),
.x2960(x2960),
.x2961(x2961),
.x2962(x2962),
.x2963(x2963),
.x2964(x2964),
.x2965(x2965),
.x2966(x2966),
.x2967(x2967),
.x2968(x2968),
.x2969(x2969),
.x2970(x2970),
.x2971(x2971),
.x2972(x2972),
.x2973(x2973),
.x2974(x2974),
.x2975(x2975),
.x2976(x2976),
.x2977(x2977),
.x2978(x2978),
.x2979(x2979),
.x2980(x2980),
.x2981(x2981),
.x2982(x2982),
.x2983(x2983),
.x2984(x2984),
.x2985(x2985),
.x2986(x2986),
.x2987(x2987),
.x2988(x2988),
.x2989(x2989),
.x2990(x2990),
.x2991(x2991),
.x2992(x2992),
.x2993(x2993),
.x2994(x2994),
.x2995(x2995),
.x2996(x2996),
.x2997(x2997),
.x2998(x2998),
.x2999(x2999),
.x3000(x3000),
.x3001(x3001),
.x3002(x3002),
.x3003(x3003),
.x3004(x3004),
.x3005(x3005),
.x3006(x3006),
.x3007(x3007),
.x3008(x3008),
.x3009(x3009),
.x3010(x3010),
.x3011(x3011),
.x3012(x3012),
.x3013(x3013),
.x3014(x3014),
.x3015(x3015),
.x3016(x3016),
.x3017(x3017),
.x3018(x3018),
.x3019(x3019),
.x3020(x3020),
.x3021(x3021),
.x3022(x3022),
.x3023(x3023),
.x3024(x3024),
.x3025(x3025),
.x3026(x3026),
.x3027(x3027),
.x3028(x3028),
.x3029(x3029),
.x3030(x3030),
.x3031(x3031),
.x3032(x3032),
.x3033(x3033),
.x3034(x3034),
.x3035(x3035),
.x3036(x3036),
.x3037(x3037),
.x3038(x3038),
.x3039(x3039),
.x3040(x3040),
.x3041(x3041),
.x3042(x3042),
.x3043(x3043),
.x3044(x3044),
.x3045(x3045),
.x3046(x3046),
.x3047(x3047),
.x3048(x3048),
.x3049(x3049),
.x3050(x3050),
.x3051(x3051),
.x3052(x3052),
.x3053(x3053),
.x3054(x3054),
.x3055(x3055),
.x3056(x3056),
.x3057(x3057),
.x3058(x3058),
.x3059(x3059),
.x3060(x3060),
.x3061(x3061),
.x3062(x3062),
.x3063(x3063),
.x3064(x3064),
.x3065(x3065),
.x3066(x3066),
.x3067(x3067),
.x3068(x3068),
.x3069(x3069),
.x3070(x3070),
.x3071(x3071),
.y0(conv11in[0]),
.y1(conv11in[1]),
.y2(conv11in[2]),
.y3(conv11in[3]),
.y4(conv11in[4]),
.y5(conv11in[5]),
.y6(conv11in[6]),
.y7(conv11in[7]),
.y8(conv11in[8]),
.y9(conv11in[9]),
.y10(conv11in[10]),
.y11(conv11in[11]),
.y12(conv11in[12]),
.y13(conv11in[13]),
.y14(conv11in[14]),
.y15(conv11in[15]),
.y16(conv11in[16]),
.y17(conv11in[17]),
.y18(conv11in[18]),
.y19(conv11in[19]),
.y20(conv11in[20]),
.y21(conv11in[21]),
.y22(conv11in[22]),
.y23(conv11in[23]),
.y24(conv11in[24]),
.y25(conv11in[25]),
.y26(conv11in[26]),
.y27(conv11in[27]),
.y28(conv11in[28]),
.y29(conv11in[29]),
.y30(conv11in[30]),
.y31(conv11in[31]),
.y32(conv11in[32]),
.y33(conv11in[33]),
.y34(conv11in[34]),
.y35(conv11in[35]),
.y36(conv11in[36]),
.y37(conv11in[37]),
.y38(conv11in[38]),
.y39(conv11in[39]),
.y40(conv11in[40]),
.y41(conv11in[41]),
.y42(conv11in[42]),
.y43(conv11in[43]),
.y44(conv11in[44]),
.y45(conv11in[45]),
.y46(conv11in[46]),
.y47(conv11in[47]),
.y48(conv11in[48]),
.y49(conv11in[49]),
.y50(conv11in[50]),
.y51(conv11in[51]),
.y52(conv11in[52]),
.y53(conv11in[53]),
.y54(conv11in[54]),
.y55(conv11in[55]),
.y56(conv11in[56]),
.y57(conv11in[57]),
.y58(conv11in[58]),
.y59(conv11in[59]),
.y60(conv11in[60]),
.y61(conv11in[61]),
.y62(conv11in[62]),
.y63(conv11in[63]),
.y64(conv11in[64]),
.y65(conv11in[65]),
.y66(conv11in[66]),
.y67(conv11in[67]),
.y68(conv11in[68]),
.y69(conv11in[69]),
.y70(conv11in[70]),
.y71(conv11in[71]),
.y72(conv11in[72]),
.y73(conv11in[73]),
.y74(conv11in[74]),
.y75(conv11in[75]),
.y76(conv11in[76]),
.y77(conv11in[77]),
.y78(conv11in[78]),
.y79(conv11in[79]),
.y80(conv11in[80]),
.y81(conv11in[81]),
.y82(conv11in[82]),
.y83(conv11in[83]),
.y84(conv11in[84]),
.y85(conv11in[85]),
.y86(conv11in[86]),
.y87(conv11in[87]),
.y88(conv11in[88]),
.y89(conv11in[89]),
.y90(conv11in[90]),
.y91(conv11in[91]),
.y92(conv11in[92]),
.y93(conv11in[93]),
.y94(conv11in[94]),
.y95(conv11in[95]),
.y96(conv11in[96]),
.y97(conv11in[97]),
.y98(conv11in[98]),
.y99(conv11in[99]),
.y100(conv11in[100]),
.y101(conv11in[101]),
.y102(conv11in[102]),
.y103(conv11in[103]),
.y104(conv11in[104]),
.y105(conv11in[105]),
.y106(conv11in[106]),
.y107(conv11in[107]),
.y108(conv11in[108]),
.y109(conv11in[109]),
.y110(conv11in[110]),
.y111(conv11in[111]),
.y112(conv11in[112]),
.y113(conv11in[113]),
.y114(conv11in[114]),
.y115(conv11in[115]),
.y116(conv11in[116]),
.y117(conv11in[117]),
.y118(conv11in[118]),
.y119(conv11in[119]),
.y120(conv11in[120]),
.y121(conv11in[121]),
.y122(conv11in[122]),
.y123(conv11in[123]),
.y124(conv11in[124]),
.y125(conv11in[125]),
.y126(conv11in[126]),
.y127(conv11in[127]),
.y128(conv11in[128]),
.y129(conv11in[129]),
.y130(conv11in[130]),
.y131(conv11in[131]),
.y132(conv11in[132]),
.y133(conv11in[133]),
.y134(conv11in[134]),
.y135(conv11in[135]),
.y136(conv11in[136]),
.y137(conv11in[137]),
.y138(conv11in[138]),
.y139(conv11in[139]),
.y140(conv11in[140]),
.y141(conv11in[141]),
.y142(conv11in[142]),
.y143(conv11in[143]),
.y144(conv11in[144]),
.y145(conv11in[145]),
.y146(conv11in[146]),
.y147(conv11in[147]),
.y148(conv11in[148]),
.y149(conv11in[149]),
.y150(conv11in[150]),
.y151(conv11in[151]),
.y152(conv11in[152]),
.y153(conv11in[153]),
.y154(conv11in[154]),
.y155(conv11in[155]),
.y156(conv11in[156]),
.y157(conv11in[157]),
.y158(conv11in[158]),
.y159(conv11in[159]),
.y160(conv11in[160]),
.y161(conv11in[161]),
.y162(conv11in[162]),
.y163(conv11in[163]),
.y164(conv11in[164]),
.y165(conv11in[165]),
.y166(conv11in[166]),
.y167(conv11in[167]),
.y168(conv11in[168]),
.y169(conv11in[169]),
.y170(conv11in[170]),
.y171(conv11in[171]),
.y172(conv11in[172]),
.y173(conv11in[173]),
.y174(conv11in[174]),
.y175(conv11in[175]),
.y176(conv11in[176]),
.y177(conv11in[177]),
.y178(conv11in[178]),
.y179(conv11in[179]),
.y180(conv11in[180]),
.y181(conv11in[181]),
.y182(conv11in[182]),
.y183(conv11in[183]),
.y184(conv11in[184]),
.y185(conv11in[185]),
.y186(conv11in[186]),
.y187(conv11in[187]),
.y188(conv11in[188]),
.y189(conv11in[189]),
.y190(conv11in[190]),
.y191(conv11in[191]),
.y192(conv11in[192]),
.y193(conv11in[193]),
.y194(conv11in[194]),
.y195(conv11in[195]),
.y196(conv11in[196]),
.y197(conv11in[197]),
.y198(conv11in[198]),
.y199(conv11in[199]),
.y200(conv11in[200]),
.y201(conv11in[201]),
.y202(conv11in[202]),
.y203(conv11in[203]),
.y204(conv11in[204]),
.y205(conv11in[205]),
.y206(conv11in[206]),
.y207(conv11in[207]),
.y208(conv11in[208]),
.y209(conv11in[209]),
.y210(conv11in[210]),
.y211(conv11in[211]),
.y212(conv11in[212]),
.y213(conv11in[213]),
.y214(conv11in[214]),
.y215(conv11in[215]),
.y216(conv11in[216]),
.y217(conv11in[217]),
.y218(conv11in[218]),
.y219(conv11in[219]),
.y220(conv11in[220]),
.y221(conv11in[221]),
.y222(conv11in[222]),
.y223(conv11in[223]),
.y224(conv11in[224]),
.y225(conv11in[225]),
.y226(conv11in[226]),
.y227(conv11in[227]),
.y228(conv11in[228]),
.y229(conv11in[229]),
.y230(conv11in[230]),
.y231(conv11in[231]),
.y232(conv11in[232]),
.y233(conv11in[233]),
.y234(conv11in[234]),
.y235(conv11in[235]),
.y236(conv11in[236]),
.y237(conv11in[237]),
.y238(conv11in[238]),
.y239(conv11in[239]),
.y240(conv11in[240]),
.y241(conv11in[241]),
.y242(conv11in[242]),
.y243(conv11in[243]),
.y244(conv11in[244]),
.y245(conv11in[245]),
.y246(conv11in[246]),
.y247(conv11in[247]),
.y248(conv11in[248]),
.y249(conv11in[249]),
.y250(conv11in[250]),
.y251(conv11in[251]),
.y252(conv11in[252]),
.y253(conv11in[253]),
.y254(conv11in[254]),
.y255(conv11in[255]),
.y256(conv11in[256]),
.y257(conv11in[257]),
.y258(conv11in[258]),
.y259(conv11in[259]),
.y260(conv11in[260]),
.y261(conv11in[261]),
.y262(conv11in[262]),
.y263(conv11in[263]),
.y264(conv11in[264]),
.y265(conv11in[265]),
.y266(conv11in[266]),
.y267(conv11in[267]),
.y268(conv11in[268]),
.y269(conv11in[269]),
.y270(conv11in[270]),
.y271(conv11in[271]),
.y272(conv11in[272]),
.y273(conv11in[273]),
.y274(conv11in[274]),
.y275(conv11in[275]),
.y276(conv11in[276]),
.y277(conv11in[277]),
.y278(conv11in[278]),
.y279(conv11in[279]),
.y280(conv11in[280]),
.y281(conv11in[281]),
.y282(conv11in[282]),
.y283(conv11in[283]),
.y284(conv11in[284]),
.y285(conv11in[285]),
.y286(conv11in[286]),
.y287(conv11in[287]),
.y288(conv11in[288]),
.y289(conv11in[289]),
.y290(conv11in[290]),
.y291(conv11in[291]),
.y292(conv11in[292]),
.y293(conv11in[293]),
.y294(conv11in[294]),
.y295(conv11in[295]),
.y296(conv11in[296]),
.y297(conv11in[297]),
.y298(conv11in[298]),
.y299(conv11in[299]),
.y300(conv11in[300]),
.y301(conv11in[301]),
.y302(conv11in[302]),
.y303(conv11in[303]),
.y304(conv11in[304]),
.y305(conv11in[305]),
.y306(conv11in[306]),
.y307(conv11in[307]),
.y308(conv11in[308]),
.y309(conv11in[309]),
.y310(conv11in[310]),
.y311(conv11in[311]),
.y312(conv11in[312]),
.y313(conv11in[313]),
.y314(conv11in[314]),
.y315(conv11in[315]),
.y316(conv11in[316]),
.y317(conv11in[317]),
.y318(conv11in[318]),
.y319(conv11in[319]),
.y320(conv11in[320]),
.y321(conv11in[321]),
.y322(conv11in[322]),
.y323(conv11in[323]),
.y324(conv11in[324]),
.y325(conv11in[325]),
.y326(conv11in[326]),
.y327(conv11in[327]),
.y328(conv11in[328]),
.y329(conv11in[329]),
.y330(conv11in[330]),
.y331(conv11in[331]),
.y332(conv11in[332]),
.y333(conv11in[333]),
.y334(conv11in[334]),
.y335(conv11in[335]),
.y336(conv11in[336]),
.y337(conv11in[337]),
.y338(conv11in[338]),
.y339(conv11in[339]),
.y340(conv11in[340]),
.y341(conv11in[341]),
.y342(conv11in[342]),
.y343(conv11in[343]),
.y344(conv11in[344]),
.y345(conv11in[345]),
.y346(conv11in[346]),
.y347(conv11in[347]),
.y348(conv11in[348]),
.y349(conv11in[349]),
.y350(conv11in[350]),
.y351(conv11in[351]),
.y352(conv11in[352]),
.y353(conv11in[353]),
.y354(conv11in[354]),
.y355(conv11in[355]),
.y356(conv11in[356]),
.y357(conv11in[357]),
.y358(conv11in[358]),
.y359(conv11in[359]),
.y360(conv11in[360]),
.y361(conv11in[361]),
.y362(conv11in[362]),
.y363(conv11in[363]),
.y364(conv11in[364]),
.y365(conv11in[365]),
.y366(conv11in[366]),
.y367(conv11in[367]),
.y368(conv11in[368]),
.y369(conv11in[369]),
.y370(conv11in[370]),
.y371(conv11in[371]),
.y372(conv11in[372]),
.y373(conv11in[373]),
.y374(conv11in[374]),
.y375(conv11in[375]),
.y376(conv11in[376]),
.y377(conv11in[377]),
.y378(conv11in[378]),
.y379(conv11in[379]),
.y380(conv11in[380]),
.y381(conv11in[381]),
.y382(conv11in[382]),
.y383(conv11in[383]),
.y384(conv11in[384]),
.y385(conv11in[385]),
.y386(conv11in[386]),
.y387(conv11in[387]),
.y388(conv11in[388]),
.y389(conv11in[389]),
.y390(conv11in[390]),
.y391(conv11in[391]),
.y392(conv11in[392]),
.y393(conv11in[393]),
.y394(conv11in[394]),
.y395(conv11in[395]),
.y396(conv11in[396]),
.y397(conv11in[397]),
.y398(conv11in[398]),
.y399(conv11in[399]),
.y400(conv11in[400]),
.y401(conv11in[401]),
.y402(conv11in[402]),
.y403(conv11in[403]),
.y404(conv11in[404]),
.y405(conv11in[405]),
.y406(conv11in[406]),
.y407(conv11in[407]),
.y408(conv11in[408]),
.y409(conv11in[409]),
.y410(conv11in[410]),
.y411(conv11in[411]),
.y412(conv11in[412]),
.y413(conv11in[413]),
.y414(conv11in[414]),
.y415(conv11in[415]),
.y416(conv11in[416]),
.y417(conv11in[417]),
.y418(conv11in[418]),
.y419(conv11in[419]),
.y420(conv11in[420]),
.y421(conv11in[421]),
.y422(conv11in[422]),
.y423(conv11in[423]),
.y424(conv11in[424]),
.y425(conv11in[425]),
.y426(conv11in[426]),
.y427(conv11in[427]),
.y428(conv11in[428]),
.y429(conv11in[429]),
.y430(conv11in[430]),
.y431(conv11in[431]),
.y432(conv11in[432]),
.y433(conv11in[433]),
.y434(conv11in[434]),
.y435(conv11in[435]),
.y436(conv11in[436]),
.y437(conv11in[437]),
.y438(conv11in[438]),
.y439(conv11in[439]),
.y440(conv11in[440]),
.y441(conv11in[441]),
.y442(conv11in[442]),
.y443(conv11in[443]),
.y444(conv11in[444]),
.y445(conv11in[445]),
.y446(conv11in[446]),
.y447(conv11in[447]),
.y448(conv11in[448]),
.y449(conv11in[449]),
.y450(conv11in[450]),
.y451(conv11in[451]),
.y452(conv11in[452]),
.y453(conv11in[453]),
.y454(conv11in[454]),
.y455(conv11in[455]),
.y456(conv11in[456]),
.y457(conv11in[457]),
.y458(conv11in[458]),
.y459(conv11in[459]),
.y460(conv11in[460]),
.y461(conv11in[461]),
.y462(conv11in[462]),
.y463(conv11in[463]),
.y464(conv11in[464]),
.y465(conv11in[465]),
.y466(conv11in[466]),
.y467(conv11in[467]),
.y468(conv11in[468]),
.y469(conv11in[469]),
.y470(conv11in[470]),
.y471(conv11in[471]),
.y472(conv11in[472]),
.y473(conv11in[473]),
.y474(conv11in[474]),
.y475(conv11in[475]),
.y476(conv11in[476]),
.y477(conv11in[477]),
.y478(conv11in[478]),
.y479(conv11in[479]),
.y480(conv11in[480]),
.y481(conv11in[481]),
.y482(conv11in[482]),
.y483(conv11in[483]),
.y484(conv11in[484]),
.y485(conv11in[485]),
.y486(conv11in[486]),
.y487(conv11in[487]),
.y488(conv11in[488]),
.y489(conv11in[489]),
.y490(conv11in[490]),
.y491(conv11in[491]),
.y492(conv11in[492]),
.y493(conv11in[493]),
.y494(conv11in[494]),
.y495(conv11in[495]),
.y496(conv11in[496]),
.y497(conv11in[497]),
.y498(conv11in[498]),
.y499(conv11in[499]),
.y500(conv11in[500]),
.y501(conv11in[501]),
.y502(conv11in[502]),
.y503(conv11in[503]),
.y504(conv11in[504]),
.y505(conv11in[505]),
.y506(conv11in[506]),
.y507(conv11in[507]),
.y508(conv11in[508]),
.y509(conv11in[509]),
.y510(conv11in[510]),
.y511(conv11in[511]),
.y512(conv11in[512]),
.y513(conv11in[513]),
.y514(conv11in[514]),
.y515(conv11in[515]),
.y516(conv11in[516]),
.y517(conv11in[517]),
.y518(conv11in[518]),
.y519(conv11in[519]),
.y520(conv11in[520]),
.y521(conv11in[521]),
.y522(conv11in[522]),
.y523(conv11in[523]),
.y524(conv11in[524]),
.y525(conv11in[525]),
.y526(conv11in[526]),
.y527(conv11in[527]),
.y528(conv11in[528]),
.y529(conv11in[529]),
.y530(conv11in[530]),
.y531(conv11in[531]),
.y532(conv11in[532]),
.y533(conv11in[533]),
.y534(conv11in[534]),
.y535(conv11in[535]),
.y536(conv11in[536]),
.y537(conv11in[537]),
.y538(conv11in[538]),
.y539(conv11in[539]),
.y540(conv11in[540]),
.y541(conv11in[541]),
.y542(conv11in[542]),
.y543(conv11in[543]),
.y544(conv11in[544]),
.y545(conv11in[545]),
.y546(conv11in[546]),
.y547(conv11in[547]),
.y548(conv11in[548]),
.y549(conv11in[549]),
.y550(conv11in[550]),
.y551(conv11in[551]),
.y552(conv11in[552]),
.y553(conv11in[553]),
.y554(conv11in[554]),
.y555(conv11in[555]),
.y556(conv11in[556]),
.y557(conv11in[557]),
.y558(conv11in[558]),
.y559(conv11in[559]),
.y560(conv11in[560]),
.y561(conv11in[561]),
.y562(conv11in[562]),
.y563(conv11in[563]),
.y564(conv11in[564]),
.y565(conv11in[565]),
.y566(conv11in[566]),
.y567(conv11in[567]),
.y568(conv11in[568]),
.y569(conv11in[569]),
.y570(conv11in[570]),
.y571(conv11in[571]),
.y572(conv11in[572]),
.y573(conv11in[573]),
.y574(conv11in[574]),
.y575(conv11in[575]),
.y576(conv11in[576]),
.y577(conv11in[577]),
.y578(conv11in[578]),
.y579(conv11in[579]),
.y580(conv11in[580]),
.y581(conv11in[581]),
.y582(conv11in[582]),
.y583(conv11in[583]),
.y584(conv11in[584]),
.y585(conv11in[585]),
.y586(conv11in[586]),
.y587(conv11in[587]),
.y588(conv11in[588]),
.y589(conv11in[589]),
.y590(conv11in[590]),
.y591(conv11in[591]),
.y592(conv11in[592]),
.y593(conv11in[593]),
.y594(conv11in[594]),
.y595(conv11in[595]),
.y596(conv11in[596]),
.y597(conv11in[597]),
.y598(conv11in[598]),
.y599(conv11in[599]),
.y600(conv11in[600]),
.y601(conv11in[601]),
.y602(conv11in[602]),
.y603(conv11in[603]),
.y604(conv11in[604]),
.y605(conv11in[605]),
.y606(conv11in[606]),
.y607(conv11in[607]),
.y608(conv11in[608]),
.y609(conv11in[609]),
.y610(conv11in[610]),
.y611(conv11in[611]),
.y612(conv11in[612]),
.y613(conv11in[613]),
.y614(conv11in[614]),
.y615(conv11in[615]),
.y616(conv11in[616]),
.y617(conv11in[617]),
.y618(conv11in[618]),
.y619(conv11in[619]),
.y620(conv11in[620]),
.y621(conv11in[621]),
.y622(conv11in[622]),
.y623(conv11in[623]),
.y624(conv11in[624]),
.y625(conv11in[625]),
.y626(conv11in[626]),
.y627(conv11in[627]),
.y628(conv11in[628]),
.y629(conv11in[629]),
.y630(conv11in[630]),
.y631(conv11in[631]),
.y632(conv11in[632]),
.y633(conv11in[633]),
.y634(conv11in[634]),
.y635(conv11in[635]),
.y636(conv11in[636]),
.y637(conv11in[637]),
.y638(conv11in[638]),
.y639(conv11in[639]),
.y640(conv11in[640]),
.y641(conv11in[641]),
.y642(conv11in[642]),
.y643(conv11in[643]),
.y644(conv11in[644]),
.y645(conv11in[645]),
.y646(conv11in[646]),
.y647(conv11in[647]),
.y648(conv11in[648]),
.y649(conv11in[649]),
.y650(conv11in[650]),
.y651(conv11in[651]),
.y652(conv11in[652]),
.y653(conv11in[653]),
.y654(conv11in[654]),
.y655(conv11in[655]),
.y656(conv11in[656]),
.y657(conv11in[657]),
.y658(conv11in[658]),
.y659(conv11in[659]),
.y660(conv11in[660]),
.y661(conv11in[661]),
.y662(conv11in[662]),
.y663(conv11in[663]),
.y664(conv11in[664]),
.y665(conv11in[665]),
.y666(conv11in[666]),
.y667(conv11in[667]),
.y668(conv11in[668]),
.y669(conv11in[669]),
.y670(conv11in[670]),
.y671(conv11in[671]),
.y672(conv11in[672]),
.y673(conv11in[673]),
.y674(conv11in[674]),
.y675(conv11in[675]),
.y676(conv11in[676]),
.y677(conv11in[677]),
.y678(conv11in[678]),
.y679(conv11in[679]),
.y680(conv11in[680]),
.y681(conv11in[681]),
.y682(conv11in[682]),
.y683(conv11in[683]),
.y684(conv11in[684]),
.y685(conv11in[685]),
.y686(conv11in[686]),
.y687(conv11in[687]),
.y688(conv11in[688]),
.y689(conv11in[689]),
.y690(conv11in[690]),
.y691(conv11in[691]),
.y692(conv11in[692]),
.y693(conv11in[693]),
.y694(conv11in[694]),
.y695(conv11in[695]),
.y696(conv11in[696]),
.y697(conv11in[697]),
.y698(conv11in[698]),
.y699(conv11in[699]),
.y700(conv11in[700]),
.y701(conv11in[701]),
.y702(conv11in[702]),
.y703(conv11in[703]),
.y704(conv11in[704]),
.y705(conv11in[705]),
.y706(conv11in[706]),
.y707(conv11in[707]),
.y708(conv11in[708]),
.y709(conv11in[709]),
.y710(conv11in[710]),
.y711(conv11in[711]),
.y712(conv11in[712]),
.y713(conv11in[713]),
.y714(conv11in[714]),
.y715(conv11in[715]),
.y716(conv11in[716]),
.y717(conv11in[717]),
.y718(conv11in[718]),
.y719(conv11in[719]),
.y720(conv11in[720]),
.y721(conv11in[721]),
.y722(conv11in[722]),
.y723(conv11in[723]),
.y724(conv11in[724]),
.y725(conv11in[725]),
.y726(conv11in[726]),
.y727(conv11in[727]),
.y728(conv11in[728]),
.y729(conv11in[729]),
.y730(conv11in[730]),
.y731(conv11in[731]),
.y732(conv11in[732]),
.y733(conv11in[733]),
.y734(conv11in[734]),
.y735(conv11in[735]),
.y736(conv11in[736]),
.y737(conv11in[737]),
.y738(conv11in[738]),
.y739(conv11in[739]),
.y740(conv11in[740]),
.y741(conv11in[741]),
.y742(conv11in[742]),
.y743(conv11in[743]),
.y744(conv11in[744]),
.y745(conv11in[745]),
.y746(conv11in[746]),
.y747(conv11in[747]),
.y748(conv11in[748]),
.y749(conv11in[749]),
.y750(conv11in[750]),
.y751(conv11in[751]),
.y752(conv11in[752]),
.y753(conv11in[753]),
.y754(conv11in[754]),
.y755(conv11in[755]),
.y756(conv11in[756]),
.y757(conv11in[757]),
.y758(conv11in[758]),
.y759(conv11in[759]),
.y760(conv11in[760]),
.y761(conv11in[761]),
.y762(conv11in[762]),
.y763(conv11in[763]),
.y764(conv11in[764]),
.y765(conv11in[765]),
.y766(conv11in[766]),
.y767(conv11in[767]) );
wire [4:0]conv11out[0:8*8*10-1];
wire [4:0]conv21out[0:4*4*18-1];
wire [4:0]conv22out[0:4*4*13-1];
wire [5:0]dense1out[0:20-1];
Conv11 conv11(.x0(conv11in[0]),
.x1(conv11in[1]),
.x2(conv11in[2]),
.x3(conv11in[3]),
.x4(conv11in[4]),
.x5(conv11in[5]),
.x6(conv11in[6]),
.x7(conv11in[7]),
.x8(conv11in[8]),
.x9(conv11in[9]),
.x10(conv11in[10]),
.x11(conv11in[11]),
.x12(conv11in[12]),
.x13(conv11in[13]),
.x14(conv11in[14]),
.x15(conv11in[15]),
.x16(conv11in[16]),
.x17(conv11in[17]),
.x18(conv11in[18]),
.x19(conv11in[19]),
.x20(conv11in[20]),
.x21(conv11in[21]),
.x22(conv11in[22]),
.x23(conv11in[23]),
.x24(conv11in[24]),
.x25(conv11in[25]),
.x26(conv11in[26]),
.x27(conv11in[27]),
.x28(conv11in[28]),
.x29(conv11in[29]),
.x30(conv11in[30]),
.x31(conv11in[31]),
.x32(conv11in[32]),
.x33(conv11in[33]),
.x34(conv11in[34]),
.x35(conv11in[35]),
.x36(conv11in[36]),
.x37(conv11in[37]),
.x38(conv11in[38]),
.x39(conv11in[39]),
.x40(conv11in[40]),
.x41(conv11in[41]),
.x42(conv11in[42]),
.x43(conv11in[43]),
.x44(conv11in[44]),
.x45(conv11in[45]),
.x46(conv11in[46]),
.x47(conv11in[47]),
.x48(conv11in[48]),
.x49(conv11in[49]),
.x50(conv11in[50]),
.x51(conv11in[51]),
.x52(conv11in[52]),
.x53(conv11in[53]),
.x54(conv11in[54]),
.x55(conv11in[55]),
.x56(conv11in[56]),
.x57(conv11in[57]),
.x58(conv11in[58]),
.x59(conv11in[59]),
.x60(conv11in[60]),
.x61(conv11in[61]),
.x62(conv11in[62]),
.x63(conv11in[63]),
.x64(conv11in[64]),
.x65(conv11in[65]),
.x66(conv11in[66]),
.x67(conv11in[67]),
.x68(conv11in[68]),
.x69(conv11in[69]),
.x70(conv11in[70]),
.x71(conv11in[71]),
.x72(conv11in[72]),
.x73(conv11in[73]),
.x74(conv11in[74]),
.x75(conv11in[75]),
.x76(conv11in[76]),
.x77(conv11in[77]),
.x78(conv11in[78]),
.x79(conv11in[79]),
.x80(conv11in[80]),
.x81(conv11in[81]),
.x82(conv11in[82]),
.x83(conv11in[83]),
.x84(conv11in[84]),
.x85(conv11in[85]),
.x86(conv11in[86]),
.x87(conv11in[87]),
.x88(conv11in[88]),
.x89(conv11in[89]),
.x90(conv11in[90]),
.x91(conv11in[91]),
.x92(conv11in[92]),
.x93(conv11in[93]),
.x94(conv11in[94]),
.x95(conv11in[95]),
.x96(conv11in[96]),
.x97(conv11in[97]),
.x98(conv11in[98]),
.x99(conv11in[99]),
.x100(conv11in[100]),
.x101(conv11in[101]),
.x102(conv11in[102]),
.x103(conv11in[103]),
.x104(conv11in[104]),
.x105(conv11in[105]),
.x106(conv11in[106]),
.x107(conv11in[107]),
.x108(conv11in[108]),
.x109(conv11in[109]),
.x110(conv11in[110]),
.x111(conv11in[111]),
.x112(conv11in[112]),
.x113(conv11in[113]),
.x114(conv11in[114]),
.x115(conv11in[115]),
.x116(conv11in[116]),
.x117(conv11in[117]),
.x118(conv11in[118]),
.x119(conv11in[119]),
.x120(conv11in[120]),
.x121(conv11in[121]),
.x122(conv11in[122]),
.x123(conv11in[123]),
.x124(conv11in[124]),
.x125(conv11in[125]),
.x126(conv11in[126]),
.x127(conv11in[127]),
.x128(conv11in[128]),
.x129(conv11in[129]),
.x130(conv11in[130]),
.x131(conv11in[131]),
.x132(conv11in[132]),
.x133(conv11in[133]),
.x134(conv11in[134]),
.x135(conv11in[135]),
.x136(conv11in[136]),
.x137(conv11in[137]),
.x138(conv11in[138]),
.x139(conv11in[139]),
.x140(conv11in[140]),
.x141(conv11in[141]),
.x142(conv11in[142]),
.x143(conv11in[143]),
.x144(conv11in[144]),
.x145(conv11in[145]),
.x146(conv11in[146]),
.x147(conv11in[147]),
.x148(conv11in[148]),
.x149(conv11in[149]),
.x150(conv11in[150]),
.x151(conv11in[151]),
.x152(conv11in[152]),
.x153(conv11in[153]),
.x154(conv11in[154]),
.x155(conv11in[155]),
.x156(conv11in[156]),
.x157(conv11in[157]),
.x158(conv11in[158]),
.x159(conv11in[159]),
.x160(conv11in[160]),
.x161(conv11in[161]),
.x162(conv11in[162]),
.x163(conv11in[163]),
.x164(conv11in[164]),
.x165(conv11in[165]),
.x166(conv11in[166]),
.x167(conv11in[167]),
.x168(conv11in[168]),
.x169(conv11in[169]),
.x170(conv11in[170]),
.x171(conv11in[171]),
.x172(conv11in[172]),
.x173(conv11in[173]),
.x174(conv11in[174]),
.x175(conv11in[175]),
.x176(conv11in[176]),
.x177(conv11in[177]),
.x178(conv11in[178]),
.x179(conv11in[179]),
.x180(conv11in[180]),
.x181(conv11in[181]),
.x182(conv11in[182]),
.x183(conv11in[183]),
.x184(conv11in[184]),
.x185(conv11in[185]),
.x186(conv11in[186]),
.x187(conv11in[187]),
.x188(conv11in[188]),
.x189(conv11in[189]),
.x190(conv11in[190]),
.x191(conv11in[191]),
.x192(conv11in[192]),
.x193(conv11in[193]),
.x194(conv11in[194]),
.x195(conv11in[195]),
.x196(conv11in[196]),
.x197(conv11in[197]),
.x198(conv11in[198]),
.x199(conv11in[199]),
.x200(conv11in[200]),
.x201(conv11in[201]),
.x202(conv11in[202]),
.x203(conv11in[203]),
.x204(conv11in[204]),
.x205(conv11in[205]),
.x206(conv11in[206]),
.x207(conv11in[207]),
.x208(conv11in[208]),
.x209(conv11in[209]),
.x210(conv11in[210]),
.x211(conv11in[211]),
.x212(conv11in[212]),
.x213(conv11in[213]),
.x214(conv11in[214]),
.x215(conv11in[215]),
.x216(conv11in[216]),
.x217(conv11in[217]),
.x218(conv11in[218]),
.x219(conv11in[219]),
.x220(conv11in[220]),
.x221(conv11in[221]),
.x222(conv11in[222]),
.x223(conv11in[223]),
.x224(conv11in[224]),
.x225(conv11in[225]),
.x226(conv11in[226]),
.x227(conv11in[227]),
.x228(conv11in[228]),
.x229(conv11in[229]),
.x230(conv11in[230]),
.x231(conv11in[231]),
.x232(conv11in[232]),
.x233(conv11in[233]),
.x234(conv11in[234]),
.x235(conv11in[235]),
.x236(conv11in[236]),
.x237(conv11in[237]),
.x238(conv11in[238]),
.x239(conv11in[239]),
.x240(conv11in[240]),
.x241(conv11in[241]),
.x242(conv11in[242]),
.x243(conv11in[243]),
.x244(conv11in[244]),
.x245(conv11in[245]),
.x246(conv11in[246]),
.x247(conv11in[247]),
.x248(conv11in[248]),
.x249(conv11in[249]),
.x250(conv11in[250]),
.x251(conv11in[251]),
.x252(conv11in[252]),
.x253(conv11in[253]),
.x254(conv11in[254]),
.x255(conv11in[255]),
.x256(conv11in[256]),
.x257(conv11in[257]),
.x258(conv11in[258]),
.x259(conv11in[259]),
.x260(conv11in[260]),
.x261(conv11in[261]),
.x262(conv11in[262]),
.x263(conv11in[263]),
.x264(conv11in[264]),
.x265(conv11in[265]),
.x266(conv11in[266]),
.x267(conv11in[267]),
.x268(conv11in[268]),
.x269(conv11in[269]),
.x270(conv11in[270]),
.x271(conv11in[271]),
.x272(conv11in[272]),
.x273(conv11in[273]),
.x274(conv11in[274]),
.x275(conv11in[275]),
.x276(conv11in[276]),
.x277(conv11in[277]),
.x278(conv11in[278]),
.x279(conv11in[279]),
.x280(conv11in[280]),
.x281(conv11in[281]),
.x282(conv11in[282]),
.x283(conv11in[283]),
.x284(conv11in[284]),
.x285(conv11in[285]),
.x286(conv11in[286]),
.x287(conv11in[287]),
.x288(conv11in[288]),
.x289(conv11in[289]),
.x290(conv11in[290]),
.x291(conv11in[291]),
.x292(conv11in[292]),
.x293(conv11in[293]),
.x294(conv11in[294]),
.x295(conv11in[295]),
.x296(conv11in[296]),
.x297(conv11in[297]),
.x298(conv11in[298]),
.x299(conv11in[299]),
.x300(conv11in[300]),
.x301(conv11in[301]),
.x302(conv11in[302]),
.x303(conv11in[303]),
.x304(conv11in[304]),
.x305(conv11in[305]),
.x306(conv11in[306]),
.x307(conv11in[307]),
.x308(conv11in[308]),
.x309(conv11in[309]),
.x310(conv11in[310]),
.x311(conv11in[311]),
.x312(conv11in[312]),
.x313(conv11in[313]),
.x314(conv11in[314]),
.x315(conv11in[315]),
.x316(conv11in[316]),
.x317(conv11in[317]),
.x318(conv11in[318]),
.x319(conv11in[319]),
.x320(conv11in[320]),
.x321(conv11in[321]),
.x322(conv11in[322]),
.x323(conv11in[323]),
.x324(conv11in[324]),
.x325(conv11in[325]),
.x326(conv11in[326]),
.x327(conv11in[327]),
.x328(conv11in[328]),
.x329(conv11in[329]),
.x330(conv11in[330]),
.x331(conv11in[331]),
.x332(conv11in[332]),
.x333(conv11in[333]),
.x334(conv11in[334]),
.x335(conv11in[335]),
.x336(conv11in[336]),
.x337(conv11in[337]),
.x338(conv11in[338]),
.x339(conv11in[339]),
.x340(conv11in[340]),
.x341(conv11in[341]),
.x342(conv11in[342]),
.x343(conv11in[343]),
.x344(conv11in[344]),
.x345(conv11in[345]),
.x346(conv11in[346]),
.x347(conv11in[347]),
.x348(conv11in[348]),
.x349(conv11in[349]),
.x350(conv11in[350]),
.x351(conv11in[351]),
.x352(conv11in[352]),
.x353(conv11in[353]),
.x354(conv11in[354]),
.x355(conv11in[355]),
.x356(conv11in[356]),
.x357(conv11in[357]),
.x358(conv11in[358]),
.x359(conv11in[359]),
.x360(conv11in[360]),
.x361(conv11in[361]),
.x362(conv11in[362]),
.x363(conv11in[363]),
.x364(conv11in[364]),
.x365(conv11in[365]),
.x366(conv11in[366]),
.x367(conv11in[367]),
.x368(conv11in[368]),
.x369(conv11in[369]),
.x370(conv11in[370]),
.x371(conv11in[371]),
.x372(conv11in[372]),
.x373(conv11in[373]),
.x374(conv11in[374]),
.x375(conv11in[375]),
.x376(conv11in[376]),
.x377(conv11in[377]),
.x378(conv11in[378]),
.x379(conv11in[379]),
.x380(conv11in[380]),
.x381(conv11in[381]),
.x382(conv11in[382]),
.x383(conv11in[383]),
.x384(conv11in[384]),
.x385(conv11in[385]),
.x386(conv11in[386]),
.x387(conv11in[387]),
.x388(conv11in[388]),
.x389(conv11in[389]),
.x390(conv11in[390]),
.x391(conv11in[391]),
.x392(conv11in[392]),
.x393(conv11in[393]),
.x394(conv11in[394]),
.x395(conv11in[395]),
.x396(conv11in[396]),
.x397(conv11in[397]),
.x398(conv11in[398]),
.x399(conv11in[399]),
.x400(conv11in[400]),
.x401(conv11in[401]),
.x402(conv11in[402]),
.x403(conv11in[403]),
.x404(conv11in[404]),
.x405(conv11in[405]),
.x406(conv11in[406]),
.x407(conv11in[407]),
.x408(conv11in[408]),
.x409(conv11in[409]),
.x410(conv11in[410]),
.x411(conv11in[411]),
.x412(conv11in[412]),
.x413(conv11in[413]),
.x414(conv11in[414]),
.x415(conv11in[415]),
.x416(conv11in[416]),
.x417(conv11in[417]),
.x418(conv11in[418]),
.x419(conv11in[419]),
.x420(conv11in[420]),
.x421(conv11in[421]),
.x422(conv11in[422]),
.x423(conv11in[423]),
.x424(conv11in[424]),
.x425(conv11in[425]),
.x426(conv11in[426]),
.x427(conv11in[427]),
.x428(conv11in[428]),
.x429(conv11in[429]),
.x430(conv11in[430]),
.x431(conv11in[431]),
.x432(conv11in[432]),
.x433(conv11in[433]),
.x434(conv11in[434]),
.x435(conv11in[435]),
.x436(conv11in[436]),
.x437(conv11in[437]),
.x438(conv11in[438]),
.x439(conv11in[439]),
.x440(conv11in[440]),
.x441(conv11in[441]),
.x442(conv11in[442]),
.x443(conv11in[443]),
.x444(conv11in[444]),
.x445(conv11in[445]),
.x446(conv11in[446]),
.x447(conv11in[447]),
.x448(conv11in[448]),
.x449(conv11in[449]),
.x450(conv11in[450]),
.x451(conv11in[451]),
.x452(conv11in[452]),
.x453(conv11in[453]),
.x454(conv11in[454]),
.x455(conv11in[455]),
.x456(conv11in[456]),
.x457(conv11in[457]),
.x458(conv11in[458]),
.x459(conv11in[459]),
.x460(conv11in[460]),
.x461(conv11in[461]),
.x462(conv11in[462]),
.x463(conv11in[463]),
.x464(conv11in[464]),
.x465(conv11in[465]),
.x466(conv11in[466]),
.x467(conv11in[467]),
.x468(conv11in[468]),
.x469(conv11in[469]),
.x470(conv11in[470]),
.x471(conv11in[471]),
.x472(conv11in[472]),
.x473(conv11in[473]),
.x474(conv11in[474]),
.x475(conv11in[475]),
.x476(conv11in[476]),
.x477(conv11in[477]),
.x478(conv11in[478]),
.x479(conv11in[479]),
.x480(conv11in[480]),
.x481(conv11in[481]),
.x482(conv11in[482]),
.x483(conv11in[483]),
.x484(conv11in[484]),
.x485(conv11in[485]),
.x486(conv11in[486]),
.x487(conv11in[487]),
.x488(conv11in[488]),
.x489(conv11in[489]),
.x490(conv11in[490]),
.x491(conv11in[491]),
.x492(conv11in[492]),
.x493(conv11in[493]),
.x494(conv11in[494]),
.x495(conv11in[495]),
.x496(conv11in[496]),
.x497(conv11in[497]),
.x498(conv11in[498]),
.x499(conv11in[499]),
.x500(conv11in[500]),
.x501(conv11in[501]),
.x502(conv11in[502]),
.x503(conv11in[503]),
.x504(conv11in[504]),
.x505(conv11in[505]),
.x506(conv11in[506]),
.x507(conv11in[507]),
.x508(conv11in[508]),
.x509(conv11in[509]),
.x510(conv11in[510]),
.x511(conv11in[511]),
.x512(conv11in[512]),
.x513(conv11in[513]),
.x514(conv11in[514]),
.x515(conv11in[515]),
.x516(conv11in[516]),
.x517(conv11in[517]),
.x518(conv11in[518]),
.x519(conv11in[519]),
.x520(conv11in[520]),
.x521(conv11in[521]),
.x522(conv11in[522]),
.x523(conv11in[523]),
.x524(conv11in[524]),
.x525(conv11in[525]),
.x526(conv11in[526]),
.x527(conv11in[527]),
.x528(conv11in[528]),
.x529(conv11in[529]),
.x530(conv11in[530]),
.x531(conv11in[531]),
.x532(conv11in[532]),
.x533(conv11in[533]),
.x534(conv11in[534]),
.x535(conv11in[535]),
.x536(conv11in[536]),
.x537(conv11in[537]),
.x538(conv11in[538]),
.x539(conv11in[539]),
.x540(conv11in[540]),
.x541(conv11in[541]),
.x542(conv11in[542]),
.x543(conv11in[543]),
.x544(conv11in[544]),
.x545(conv11in[545]),
.x546(conv11in[546]),
.x547(conv11in[547]),
.x548(conv11in[548]),
.x549(conv11in[549]),
.x550(conv11in[550]),
.x551(conv11in[551]),
.x552(conv11in[552]),
.x553(conv11in[553]),
.x554(conv11in[554]),
.x555(conv11in[555]),
.x556(conv11in[556]),
.x557(conv11in[557]),
.x558(conv11in[558]),
.x559(conv11in[559]),
.x560(conv11in[560]),
.x561(conv11in[561]),
.x562(conv11in[562]),
.x563(conv11in[563]),
.x564(conv11in[564]),
.x565(conv11in[565]),
.x566(conv11in[566]),
.x567(conv11in[567]),
.x568(conv11in[568]),
.x569(conv11in[569]),
.x570(conv11in[570]),
.x571(conv11in[571]),
.x572(conv11in[572]),
.x573(conv11in[573]),
.x574(conv11in[574]),
.x575(conv11in[575]),
.x576(conv11in[576]),
.x577(conv11in[577]),
.x578(conv11in[578]),
.x579(conv11in[579]),
.x580(conv11in[580]),
.x581(conv11in[581]),
.x582(conv11in[582]),
.x583(conv11in[583]),
.x584(conv11in[584]),
.x585(conv11in[585]),
.x586(conv11in[586]),
.x587(conv11in[587]),
.x588(conv11in[588]),
.x589(conv11in[589]),
.x590(conv11in[590]),
.x591(conv11in[591]),
.x592(conv11in[592]),
.x593(conv11in[593]),
.x594(conv11in[594]),
.x595(conv11in[595]),
.x596(conv11in[596]),
.x597(conv11in[597]),
.x598(conv11in[598]),
.x599(conv11in[599]),
.x600(conv11in[600]),
.x601(conv11in[601]),
.x602(conv11in[602]),
.x603(conv11in[603]),
.x604(conv11in[604]),
.x605(conv11in[605]),
.x606(conv11in[606]),
.x607(conv11in[607]),
.x608(conv11in[608]),
.x609(conv11in[609]),
.x610(conv11in[610]),
.x611(conv11in[611]),
.x612(conv11in[612]),
.x613(conv11in[613]),
.x614(conv11in[614]),
.x615(conv11in[615]),
.x616(conv11in[616]),
.x617(conv11in[617]),
.x618(conv11in[618]),
.x619(conv11in[619]),
.x620(conv11in[620]),
.x621(conv11in[621]),
.x622(conv11in[622]),
.x623(conv11in[623]),
.x624(conv11in[624]),
.x625(conv11in[625]),
.x626(conv11in[626]),
.x627(conv11in[627]),
.x628(conv11in[628]),
.x629(conv11in[629]),
.x630(conv11in[630]),
.x631(conv11in[631]),
.x632(conv11in[632]),
.x633(conv11in[633]),
.x634(conv11in[634]),
.x635(conv11in[635]),
.x636(conv11in[636]),
.x637(conv11in[637]),
.x638(conv11in[638]),
.x639(conv11in[639]),
.x640(conv11in[640]),
.x641(conv11in[641]),
.x642(conv11in[642]),
.x643(conv11in[643]),
.x644(conv11in[644]),
.x645(conv11in[645]),
.x646(conv11in[646]),
.x647(conv11in[647]),
.x648(conv11in[648]),
.x649(conv11in[649]),
.x650(conv11in[650]),
.x651(conv11in[651]),
.x652(conv11in[652]),
.x653(conv11in[653]),
.x654(conv11in[654]),
.x655(conv11in[655]),
.x656(conv11in[656]),
.x657(conv11in[657]),
.x658(conv11in[658]),
.x659(conv11in[659]),
.x660(conv11in[660]),
.x661(conv11in[661]),
.x662(conv11in[662]),
.x663(conv11in[663]),
.x664(conv11in[664]),
.x665(conv11in[665]),
.x666(conv11in[666]),
.x667(conv11in[667]),
.x668(conv11in[668]),
.x669(conv11in[669]),
.x670(conv11in[670]),
.x671(conv11in[671]),
.x672(conv11in[672]),
.x673(conv11in[673]),
.x674(conv11in[674]),
.x675(conv11in[675]),
.x676(conv11in[676]),
.x677(conv11in[677]),
.x678(conv11in[678]),
.x679(conv11in[679]),
.x680(conv11in[680]),
.x681(conv11in[681]),
.x682(conv11in[682]),
.x683(conv11in[683]),
.x684(conv11in[684]),
.x685(conv11in[685]),
.x686(conv11in[686]),
.x687(conv11in[687]),
.x688(conv11in[688]),
.x689(conv11in[689]),
.x690(conv11in[690]),
.x691(conv11in[691]),
.x692(conv11in[692]),
.x693(conv11in[693]),
.x694(conv11in[694]),
.x695(conv11in[695]),
.x696(conv11in[696]),
.x697(conv11in[697]),
.x698(conv11in[698]),
.x699(conv11in[699]),
.x700(conv11in[700]),
.x701(conv11in[701]),
.x702(conv11in[702]),
.x703(conv11in[703]),
.x704(conv11in[704]),
.x705(conv11in[705]),
.x706(conv11in[706]),
.x707(conv11in[707]),
.x708(conv11in[708]),
.x709(conv11in[709]),
.x710(conv11in[710]),
.x711(conv11in[711]),
.x712(conv11in[712]),
.x713(conv11in[713]),
.x714(conv11in[714]),
.x715(conv11in[715]),
.x716(conv11in[716]),
.x717(conv11in[717]),
.x718(conv11in[718]),
.x719(conv11in[719]),
.x720(conv11in[720]),
.x721(conv11in[721]),
.x722(conv11in[722]),
.x723(conv11in[723]),
.x724(conv11in[724]),
.x725(conv11in[725]),
.x726(conv11in[726]),
.x727(conv11in[727]),
.x728(conv11in[728]),
.x729(conv11in[729]),
.x730(conv11in[730]),
.x731(conv11in[731]),
.x732(conv11in[732]),
.x733(conv11in[733]),
.x734(conv11in[734]),
.x735(conv11in[735]),
.x736(conv11in[736]),
.x737(conv11in[737]),
.x738(conv11in[738]),
.x739(conv11in[739]),
.x740(conv11in[740]),
.x741(conv11in[741]),
.x742(conv11in[742]),
.x743(conv11in[743]),
.x744(conv11in[744]),
.x745(conv11in[745]),
.x746(conv11in[746]),
.x747(conv11in[747]),
.x748(conv11in[748]),
.x749(conv11in[749]),
.x750(conv11in[750]),
.x751(conv11in[751]),
.x752(conv11in[752]),
.x753(conv11in[753]),
.x754(conv11in[754]),
.x755(conv11in[755]),
.x756(conv11in[756]),
.x757(conv11in[757]),
.x758(conv11in[758]),
.x759(conv11in[759]),
.x760(conv11in[760]),
.x761(conv11in[761]),
.x762(conv11in[762]),
.x763(conv11in[763]),
.x764(conv11in[764]),
.x765(conv11in[765]),
.x766(conv11in[766]),
.x767(conv11in[767]),
.y0(conv11out[0]),
.y1(conv11out[1]),
.y2(conv11out[2]),
.y3(conv11out[3]),
.y4(conv11out[4]),
.y5(conv11out[5]),
.y6(conv11out[6]),
.y7(conv11out[7]),
.y8(conv11out[8]),
.y9(conv11out[9]),
.y10(conv11out[10]),
.y11(conv11out[11]),
.y12(conv11out[12]),
.y13(conv11out[13]),
.y14(conv11out[14]),
.y15(conv11out[15]),
.y16(conv11out[16]),
.y17(conv11out[17]),
.y18(conv11out[18]),
.y19(conv11out[19]),
.y20(conv11out[20]),
.y21(conv11out[21]),
.y22(conv11out[22]),
.y23(conv11out[23]),
.y24(conv11out[24]),
.y25(conv11out[25]),
.y26(conv11out[26]),
.y27(conv11out[27]),
.y28(conv11out[28]),
.y29(conv11out[29]),
.y30(conv11out[30]),
.y31(conv11out[31]),
.y32(conv11out[32]),
.y33(conv11out[33]),
.y34(conv11out[34]),
.y35(conv11out[35]),
.y36(conv11out[36]),
.y37(conv11out[37]),
.y38(conv11out[38]),
.y39(conv11out[39]),
.y40(conv11out[40]),
.y41(conv11out[41]),
.y42(conv11out[42]),
.y43(conv11out[43]),
.y44(conv11out[44]),
.y45(conv11out[45]),
.y46(conv11out[46]),
.y47(conv11out[47]),
.y48(conv11out[48]),
.y49(conv11out[49]),
.y50(conv11out[50]),
.y51(conv11out[51]),
.y52(conv11out[52]),
.y53(conv11out[53]),
.y54(conv11out[54]),
.y55(conv11out[55]),
.y56(conv11out[56]),
.y57(conv11out[57]),
.y58(conv11out[58]),
.y59(conv11out[59]),
.y60(conv11out[60]),
.y61(conv11out[61]),
.y62(conv11out[62]),
.y63(conv11out[63]),
.y64(conv11out[64]),
.y65(conv11out[65]),
.y66(conv11out[66]),
.y67(conv11out[67]),
.y68(conv11out[68]),
.y69(conv11out[69]),
.y70(conv11out[70]),
.y71(conv11out[71]),
.y72(conv11out[72]),
.y73(conv11out[73]),
.y74(conv11out[74]),
.y75(conv11out[75]),
.y76(conv11out[76]),
.y77(conv11out[77]),
.y78(conv11out[78]),
.y79(conv11out[79]),
.y80(conv11out[80]),
.y81(conv11out[81]),
.y82(conv11out[82]),
.y83(conv11out[83]),
.y84(conv11out[84]),
.y85(conv11out[85]),
.y86(conv11out[86]),
.y87(conv11out[87]),
.y88(conv11out[88]),
.y89(conv11out[89]),
.y90(conv11out[90]),
.y91(conv11out[91]),
.y92(conv11out[92]),
.y93(conv11out[93]),
.y94(conv11out[94]),
.y95(conv11out[95]),
.y96(conv11out[96]),
.y97(conv11out[97]),
.y98(conv11out[98]),
.y99(conv11out[99]),
.y100(conv11out[100]),
.y101(conv11out[101]),
.y102(conv11out[102]),
.y103(conv11out[103]),
.y104(conv11out[104]),
.y105(conv11out[105]),
.y106(conv11out[106]),
.y107(conv11out[107]),
.y108(conv11out[108]),
.y109(conv11out[109]),
.y110(conv11out[110]),
.y111(conv11out[111]),
.y112(conv11out[112]),
.y113(conv11out[113]),
.y114(conv11out[114]),
.y115(conv11out[115]),
.y116(conv11out[116]),
.y117(conv11out[117]),
.y118(conv11out[118]),
.y119(conv11out[119]),
.y120(conv11out[120]),
.y121(conv11out[121]),
.y122(conv11out[122]),
.y123(conv11out[123]),
.y124(conv11out[124]),
.y125(conv11out[125]),
.y126(conv11out[126]),
.y127(conv11out[127]),
.y128(conv11out[128]),
.y129(conv11out[129]),
.y130(conv11out[130]),
.y131(conv11out[131]),
.y132(conv11out[132]),
.y133(conv11out[133]),
.y134(conv11out[134]),
.y135(conv11out[135]),
.y136(conv11out[136]),
.y137(conv11out[137]),
.y138(conv11out[138]),
.y139(conv11out[139]),
.y140(conv11out[140]),
.y141(conv11out[141]),
.y142(conv11out[142]),
.y143(conv11out[143]),
.y144(conv11out[144]),
.y145(conv11out[145]),
.y146(conv11out[146]),
.y147(conv11out[147]),
.y148(conv11out[148]),
.y149(conv11out[149]),
.y150(conv11out[150]),
.y151(conv11out[151]),
.y152(conv11out[152]),
.y153(conv11out[153]),
.y154(conv11out[154]),
.y155(conv11out[155]),
.y156(conv11out[156]),
.y157(conv11out[157]),
.y158(conv11out[158]),
.y159(conv11out[159]),
.y160(conv11out[160]),
.y161(conv11out[161]),
.y162(conv11out[162]),
.y163(conv11out[163]),
.y164(conv11out[164]),
.y165(conv11out[165]),
.y166(conv11out[166]),
.y167(conv11out[167]),
.y168(conv11out[168]),
.y169(conv11out[169]),
.y170(conv11out[170]),
.y171(conv11out[171]),
.y172(conv11out[172]),
.y173(conv11out[173]),
.y174(conv11out[174]),
.y175(conv11out[175]),
.y176(conv11out[176]),
.y177(conv11out[177]),
.y178(conv11out[178]),
.y179(conv11out[179]),
.y180(conv11out[180]),
.y181(conv11out[181]),
.y182(conv11out[182]),
.y183(conv11out[183]),
.y184(conv11out[184]),
.y185(conv11out[185]),
.y186(conv11out[186]),
.y187(conv11out[187]),
.y188(conv11out[188]),
.y189(conv11out[189]),
.y190(conv11out[190]),
.y191(conv11out[191]),
.y192(conv11out[192]),
.y193(conv11out[193]),
.y194(conv11out[194]),
.y195(conv11out[195]),
.y196(conv11out[196]),
.y197(conv11out[197]),
.y198(conv11out[198]),
.y199(conv11out[199]),
.y200(conv11out[200]),
.y201(conv11out[201]),
.y202(conv11out[202]),
.y203(conv11out[203]),
.y204(conv11out[204]),
.y205(conv11out[205]),
.y206(conv11out[206]),
.y207(conv11out[207]),
.y208(conv11out[208]),
.y209(conv11out[209]),
.y210(conv11out[210]),
.y211(conv11out[211]),
.y212(conv11out[212]),
.y213(conv11out[213]),
.y214(conv11out[214]),
.y215(conv11out[215]),
.y216(conv11out[216]),
.y217(conv11out[217]),
.y218(conv11out[218]),
.y219(conv11out[219]),
.y220(conv11out[220]),
.y221(conv11out[221]),
.y222(conv11out[222]),
.y223(conv11out[223]),
.y224(conv11out[224]),
.y225(conv11out[225]),
.y226(conv11out[226]),
.y227(conv11out[227]),
.y228(conv11out[228]),
.y229(conv11out[229]),
.y230(conv11out[230]),
.y231(conv11out[231]),
.y232(conv11out[232]),
.y233(conv11out[233]),
.y234(conv11out[234]),
.y235(conv11out[235]),
.y236(conv11out[236]),
.y237(conv11out[237]),
.y238(conv11out[238]),
.y239(conv11out[239]),
.y240(conv11out[240]),
.y241(conv11out[241]),
.y242(conv11out[242]),
.y243(conv11out[243]),
.y244(conv11out[244]),
.y245(conv11out[245]),
.y246(conv11out[246]),
.y247(conv11out[247]),
.y248(conv11out[248]),
.y249(conv11out[249]),
.y250(conv11out[250]),
.y251(conv11out[251]),
.y252(conv11out[252]),
.y253(conv11out[253]),
.y254(conv11out[254]),
.y255(conv11out[255]),
.y256(conv11out[256]),
.y257(conv11out[257]),
.y258(conv11out[258]),
.y259(conv11out[259]),
.y260(conv11out[260]),
.y261(conv11out[261]),
.y262(conv11out[262]),
.y263(conv11out[263]),
.y264(conv11out[264]),
.y265(conv11out[265]),
.y266(conv11out[266]),
.y267(conv11out[267]),
.y268(conv11out[268]),
.y269(conv11out[269]),
.y270(conv11out[270]),
.y271(conv11out[271]),
.y272(conv11out[272]),
.y273(conv11out[273]),
.y274(conv11out[274]),
.y275(conv11out[275]),
.y276(conv11out[276]),
.y277(conv11out[277]),
.y278(conv11out[278]),
.y279(conv11out[279]),
.y280(conv11out[280]),
.y281(conv11out[281]),
.y282(conv11out[282]),
.y283(conv11out[283]),
.y284(conv11out[284]),
.y285(conv11out[285]),
.y286(conv11out[286]),
.y287(conv11out[287]),
.y288(conv11out[288]),
.y289(conv11out[289]),
.y290(conv11out[290]),
.y291(conv11out[291]),
.y292(conv11out[292]),
.y293(conv11out[293]),
.y294(conv11out[294]),
.y295(conv11out[295]),
.y296(conv11out[296]),
.y297(conv11out[297]),
.y298(conv11out[298]),
.y299(conv11out[299]),
.y300(conv11out[300]),
.y301(conv11out[301]),
.y302(conv11out[302]),
.y303(conv11out[303]),
.y304(conv11out[304]),
.y305(conv11out[305]),
.y306(conv11out[306]),
.y307(conv11out[307]),
.y308(conv11out[308]),
.y309(conv11out[309]),
.y310(conv11out[310]),
.y311(conv11out[311]),
.y312(conv11out[312]),
.y313(conv11out[313]),
.y314(conv11out[314]),
.y315(conv11out[315]),
.y316(conv11out[316]),
.y317(conv11out[317]),
.y318(conv11out[318]),
.y319(conv11out[319]),
.y320(conv11out[320]),
.y321(conv11out[321]),
.y322(conv11out[322]),
.y323(conv11out[323]),
.y324(conv11out[324]),
.y325(conv11out[325]),
.y326(conv11out[326]),
.y327(conv11out[327]),
.y328(conv11out[328]),
.y329(conv11out[329]),
.y330(conv11out[330]),
.y331(conv11out[331]),
.y332(conv11out[332]),
.y333(conv11out[333]),
.y334(conv11out[334]),
.y335(conv11out[335]),
.y336(conv11out[336]),
.y337(conv11out[337]),
.y338(conv11out[338]),
.y339(conv11out[339]),
.y340(conv11out[340]),
.y341(conv11out[341]),
.y342(conv11out[342]),
.y343(conv11out[343]),
.y344(conv11out[344]),
.y345(conv11out[345]),
.y346(conv11out[346]),
.y347(conv11out[347]),
.y348(conv11out[348]),
.y349(conv11out[349]),
.y350(conv11out[350]),
.y351(conv11out[351]),
.y352(conv11out[352]),
.y353(conv11out[353]),
.y354(conv11out[354]),
.y355(conv11out[355]),
.y356(conv11out[356]),
.y357(conv11out[357]),
.y358(conv11out[358]),
.y359(conv11out[359]),
.y360(conv11out[360]),
.y361(conv11out[361]),
.y362(conv11out[362]),
.y363(conv11out[363]),
.y364(conv11out[364]),
.y365(conv11out[365]),
.y366(conv11out[366]),
.y367(conv11out[367]),
.y368(conv11out[368]),
.y369(conv11out[369]),
.y370(conv11out[370]),
.y371(conv11out[371]),
.y372(conv11out[372]),
.y373(conv11out[373]),
.y374(conv11out[374]),
.y375(conv11out[375]),
.y376(conv11out[376]),
.y377(conv11out[377]),
.y378(conv11out[378]),
.y379(conv11out[379]),
.y380(conv11out[380]),
.y381(conv11out[381]),
.y382(conv11out[382]),
.y383(conv11out[383]),
.y384(conv11out[384]),
.y385(conv11out[385]),
.y386(conv11out[386]),
.y387(conv11out[387]),
.y388(conv11out[388]),
.y389(conv11out[389]),
.y390(conv11out[390]),
.y391(conv11out[391]),
.y392(conv11out[392]),
.y393(conv11out[393]),
.y394(conv11out[394]),
.y395(conv11out[395]),
.y396(conv11out[396]),
.y397(conv11out[397]),
.y398(conv11out[398]),
.y399(conv11out[399]),
.y400(conv11out[400]),
.y401(conv11out[401]),
.y402(conv11out[402]),
.y403(conv11out[403]),
.y404(conv11out[404]),
.y405(conv11out[405]),
.y406(conv11out[406]),
.y407(conv11out[407]),
.y408(conv11out[408]),
.y409(conv11out[409]),
.y410(conv11out[410]),
.y411(conv11out[411]),
.y412(conv11out[412]),
.y413(conv11out[413]),
.y414(conv11out[414]),
.y415(conv11out[415]),
.y416(conv11out[416]),
.y417(conv11out[417]),
.y418(conv11out[418]),
.y419(conv11out[419]),
.y420(conv11out[420]),
.y421(conv11out[421]),
.y422(conv11out[422]),
.y423(conv11out[423]),
.y424(conv11out[424]),
.y425(conv11out[425]),
.y426(conv11out[426]),
.y427(conv11out[427]),
.y428(conv11out[428]),
.y429(conv11out[429]),
.y430(conv11out[430]),
.y431(conv11out[431]),
.y432(conv11out[432]),
.y433(conv11out[433]),
.y434(conv11out[434]),
.y435(conv11out[435]),
.y436(conv11out[436]),
.y437(conv11out[437]),
.y438(conv11out[438]),
.y439(conv11out[439]),
.y440(conv11out[440]),
.y441(conv11out[441]),
.y442(conv11out[442]),
.y443(conv11out[443]),
.y444(conv11out[444]),
.y445(conv11out[445]),
.y446(conv11out[446]),
.y447(conv11out[447]),
.y448(conv11out[448]),
.y449(conv11out[449]),
.y450(conv11out[450]),
.y451(conv11out[451]),
.y452(conv11out[452]),
.y453(conv11out[453]),
.y454(conv11out[454]),
.y455(conv11out[455]),
.y456(conv11out[456]),
.y457(conv11out[457]),
.y458(conv11out[458]),
.y459(conv11out[459]),
.y460(conv11out[460]),
.y461(conv11out[461]),
.y462(conv11out[462]),
.y463(conv11out[463]),
.y464(conv11out[464]),
.y465(conv11out[465]),
.y466(conv11out[466]),
.y467(conv11out[467]),
.y468(conv11out[468]),
.y469(conv11out[469]),
.y470(conv11out[470]),
.y471(conv11out[471]),
.y472(conv11out[472]),
.y473(conv11out[473]),
.y474(conv11out[474]),
.y475(conv11out[475]),
.y476(conv11out[476]),
.y477(conv11out[477]),
.y478(conv11out[478]),
.y479(conv11out[479]),
.y480(conv11out[480]),
.y481(conv11out[481]),
.y482(conv11out[482]),
.y483(conv11out[483]),
.y484(conv11out[484]),
.y485(conv11out[485]),
.y486(conv11out[486]),
.y487(conv11out[487]),
.y488(conv11out[488]),
.y489(conv11out[489]),
.y490(conv11out[490]),
.y491(conv11out[491]),
.y492(conv11out[492]),
.y493(conv11out[493]),
.y494(conv11out[494]),
.y495(conv11out[495]),
.y496(conv11out[496]),
.y497(conv11out[497]),
.y498(conv11out[498]),
.y499(conv11out[499]),
.y500(conv11out[500]),
.y501(conv11out[501]),
.y502(conv11out[502]),
.y503(conv11out[503]),
.y504(conv11out[504]),
.y505(conv11out[505]),
.y506(conv11out[506]),
.y507(conv11out[507]),
.y508(conv11out[508]),
.y509(conv11out[509]),
.y510(conv11out[510]),
.y511(conv11out[511]),
.y512(conv11out[512]),
.y513(conv11out[513]),
.y514(conv11out[514]),
.y515(conv11out[515]),
.y516(conv11out[516]),
.y517(conv11out[517]),
.y518(conv11out[518]),
.y519(conv11out[519]),
.y520(conv11out[520]),
.y521(conv11out[521]),
.y522(conv11out[522]),
.y523(conv11out[523]),
.y524(conv11out[524]),
.y525(conv11out[525]),
.y526(conv11out[526]),
.y527(conv11out[527]),
.y528(conv11out[528]),
.y529(conv11out[529]),
.y530(conv11out[530]),
.y531(conv11out[531]),
.y532(conv11out[532]),
.y533(conv11out[533]),
.y534(conv11out[534]),
.y535(conv11out[535]),
.y536(conv11out[536]),
.y537(conv11out[537]),
.y538(conv11out[538]),
.y539(conv11out[539]),
.y540(conv11out[540]),
.y541(conv11out[541]),
.y542(conv11out[542]),
.y543(conv11out[543]),
.y544(conv11out[544]),
.y545(conv11out[545]),
.y546(conv11out[546]),
.y547(conv11out[547]),
.y548(conv11out[548]),
.y549(conv11out[549]),
.y550(conv11out[550]),
.y551(conv11out[551]),
.y552(conv11out[552]),
.y553(conv11out[553]),
.y554(conv11out[554]),
.y555(conv11out[555]),
.y556(conv11out[556]),
.y557(conv11out[557]),
.y558(conv11out[558]),
.y559(conv11out[559]),
.y560(conv11out[560]),
.y561(conv11out[561]),
.y562(conv11out[562]),
.y563(conv11out[563]),
.y564(conv11out[564]),
.y565(conv11out[565]),
.y566(conv11out[566]),
.y567(conv11out[567]),
.y568(conv11out[568]),
.y569(conv11out[569]),
.y570(conv11out[570]),
.y571(conv11out[571]),
.y572(conv11out[572]),
.y573(conv11out[573]),
.y574(conv11out[574]),
.y575(conv11out[575]),
.y576(conv11out[576]),
.y577(conv11out[577]),
.y578(conv11out[578]),
.y579(conv11out[579]),
.y580(conv11out[580]),
.y581(conv11out[581]),
.y582(conv11out[582]),
.y583(conv11out[583]),
.y584(conv11out[584]),
.y585(conv11out[585]),
.y586(conv11out[586]),
.y587(conv11out[587]),
.y588(conv11out[588]),
.y589(conv11out[589]),
.y590(conv11out[590]),
.y591(conv11out[591]),
.y592(conv11out[592]),
.y593(conv11out[593]),
.y594(conv11out[594]),
.y595(conv11out[595]),
.y596(conv11out[596]),
.y597(conv11out[597]),
.y598(conv11out[598]),
.y599(conv11out[599]),
.y600(conv11out[600]),
.y601(conv11out[601]),
.y602(conv11out[602]),
.y603(conv11out[603]),
.y604(conv11out[604]),
.y605(conv11out[605]),
.y606(conv11out[606]),
.y607(conv11out[607]),
.y608(conv11out[608]),
.y609(conv11out[609]),
.y610(conv11out[610]),
.y611(conv11out[611]),
.y612(conv11out[612]),
.y613(conv11out[613]),
.y614(conv11out[614]),
.y615(conv11out[615]),
.y616(conv11out[616]),
.y617(conv11out[617]),
.y618(conv11out[618]),
.y619(conv11out[619]),
.y620(conv11out[620]),
.y621(conv11out[621]),
.y622(conv11out[622]),
.y623(conv11out[623]),
.y624(conv11out[624]),
.y625(conv11out[625]),
.y626(conv11out[626]),
.y627(conv11out[627]),
.y628(conv11out[628]),
.y629(conv11out[629]),
.y630(conv11out[630]),
.y631(conv11out[631]),
.y632(conv11out[632]),
.y633(conv11out[633]),
.y634(conv11out[634]),
.y635(conv11out[635]),
.y636(conv11out[636]),
.y637(conv11out[637]),
.y638(conv11out[638]),
.y639(conv11out[639]) );
Conv21 conv21(.x0(conv11out[0]),
.x1(conv11out[1]),
.x2(conv11out[2]),
.x3(conv11out[3]),
.x4(conv11out[4]),
.x5(conv11out[5]),
.x6(conv11out[6]),
.x7(conv11out[7]),
.x8(conv11out[8]),
.x9(conv11out[9]),
.x10(conv11out[10]),
.x11(conv11out[11]),
.x12(conv11out[12]),
.x13(conv11out[13]),
.x14(conv11out[14]),
.x15(conv11out[15]),
.x16(conv11out[16]),
.x17(conv11out[17]),
.x18(conv11out[18]),
.x19(conv11out[19]),
.x20(conv11out[20]),
.x21(conv11out[21]),
.x22(conv11out[22]),
.x23(conv11out[23]),
.x24(conv11out[24]),
.x25(conv11out[25]),
.x26(conv11out[26]),
.x27(conv11out[27]),
.x28(conv11out[28]),
.x29(conv11out[29]),
.x30(conv11out[30]),
.x31(conv11out[31]),
.x32(conv11out[32]),
.x33(conv11out[33]),
.x34(conv11out[34]),
.x35(conv11out[35]),
.x36(conv11out[36]),
.x37(conv11out[37]),
.x38(conv11out[38]),
.x39(conv11out[39]),
.x40(conv11out[40]),
.x41(conv11out[41]),
.x42(conv11out[42]),
.x43(conv11out[43]),
.x44(conv11out[44]),
.x45(conv11out[45]),
.x46(conv11out[46]),
.x47(conv11out[47]),
.x48(conv11out[48]),
.x49(conv11out[49]),
.x50(conv11out[50]),
.x51(conv11out[51]),
.x52(conv11out[52]),
.x53(conv11out[53]),
.x54(conv11out[54]),
.x55(conv11out[55]),
.x56(conv11out[56]),
.x57(conv11out[57]),
.x58(conv11out[58]),
.x59(conv11out[59]),
.x60(conv11out[60]),
.x61(conv11out[61]),
.x62(conv11out[62]),
.x63(conv11out[63]),
.x64(conv11out[64]),
.x65(conv11out[65]),
.x66(conv11out[66]),
.x67(conv11out[67]),
.x68(conv11out[68]),
.x69(conv11out[69]),
.x70(conv11out[70]),
.x71(conv11out[71]),
.x72(conv11out[72]),
.x73(conv11out[73]),
.x74(conv11out[74]),
.x75(conv11out[75]),
.x76(conv11out[76]),
.x77(conv11out[77]),
.x78(conv11out[78]),
.x79(conv11out[79]),
.x80(conv11out[80]),
.x81(conv11out[81]),
.x82(conv11out[82]),
.x83(conv11out[83]),
.x84(conv11out[84]),
.x85(conv11out[85]),
.x86(conv11out[86]),
.x87(conv11out[87]),
.x88(conv11out[88]),
.x89(conv11out[89]),
.x90(conv11out[90]),
.x91(conv11out[91]),
.x92(conv11out[92]),
.x93(conv11out[93]),
.x94(conv11out[94]),
.x95(conv11out[95]),
.x96(conv11out[96]),
.x97(conv11out[97]),
.x98(conv11out[98]),
.x99(conv11out[99]),
.x100(conv11out[100]),
.x101(conv11out[101]),
.x102(conv11out[102]),
.x103(conv11out[103]),
.x104(conv11out[104]),
.x105(conv11out[105]),
.x106(conv11out[106]),
.x107(conv11out[107]),
.x108(conv11out[108]),
.x109(conv11out[109]),
.x110(conv11out[110]),
.x111(conv11out[111]),
.x112(conv11out[112]),
.x113(conv11out[113]),
.x114(conv11out[114]),
.x115(conv11out[115]),
.x116(conv11out[116]),
.x117(conv11out[117]),
.x118(conv11out[118]),
.x119(conv11out[119]),
.x120(conv11out[120]),
.x121(conv11out[121]),
.x122(conv11out[122]),
.x123(conv11out[123]),
.x124(conv11out[124]),
.x125(conv11out[125]),
.x126(conv11out[126]),
.x127(conv11out[127]),
.x128(conv11out[128]),
.x129(conv11out[129]),
.x130(conv11out[130]),
.x131(conv11out[131]),
.x132(conv11out[132]),
.x133(conv11out[133]),
.x134(conv11out[134]),
.x135(conv11out[135]),
.x136(conv11out[136]),
.x137(conv11out[137]),
.x138(conv11out[138]),
.x139(conv11out[139]),
.x140(conv11out[140]),
.x141(conv11out[141]),
.x142(conv11out[142]),
.x143(conv11out[143]),
.x144(conv11out[144]),
.x145(conv11out[145]),
.x146(conv11out[146]),
.x147(conv11out[147]),
.x148(conv11out[148]),
.x149(conv11out[149]),
.x150(conv11out[150]),
.x151(conv11out[151]),
.x152(conv11out[152]),
.x153(conv11out[153]),
.x154(conv11out[154]),
.x155(conv11out[155]),
.x156(conv11out[156]),
.x157(conv11out[157]),
.x158(conv11out[158]),
.x159(conv11out[159]),
.x160(conv11out[160]),
.x161(conv11out[161]),
.x162(conv11out[162]),
.x163(conv11out[163]),
.x164(conv11out[164]),
.x165(conv11out[165]),
.x166(conv11out[166]),
.x167(conv11out[167]),
.x168(conv11out[168]),
.x169(conv11out[169]),
.x170(conv11out[170]),
.x171(conv11out[171]),
.x172(conv11out[172]),
.x173(conv11out[173]),
.x174(conv11out[174]),
.x175(conv11out[175]),
.x176(conv11out[176]),
.x177(conv11out[177]),
.x178(conv11out[178]),
.x179(conv11out[179]),
.x180(conv11out[180]),
.x181(conv11out[181]),
.x182(conv11out[182]),
.x183(conv11out[183]),
.x184(conv11out[184]),
.x185(conv11out[185]),
.x186(conv11out[186]),
.x187(conv11out[187]),
.x188(conv11out[188]),
.x189(conv11out[189]),
.x190(conv11out[190]),
.x191(conv11out[191]),
.x192(conv11out[192]),
.x193(conv11out[193]),
.x194(conv11out[194]),
.x195(conv11out[195]),
.x196(conv11out[196]),
.x197(conv11out[197]),
.x198(conv11out[198]),
.x199(conv11out[199]),
.x200(conv11out[200]),
.x201(conv11out[201]),
.x202(conv11out[202]),
.x203(conv11out[203]),
.x204(conv11out[204]),
.x205(conv11out[205]),
.x206(conv11out[206]),
.x207(conv11out[207]),
.x208(conv11out[208]),
.x209(conv11out[209]),
.x210(conv11out[210]),
.x211(conv11out[211]),
.x212(conv11out[212]),
.x213(conv11out[213]),
.x214(conv11out[214]),
.x215(conv11out[215]),
.x216(conv11out[216]),
.x217(conv11out[217]),
.x218(conv11out[218]),
.x219(conv11out[219]),
.x220(conv11out[220]),
.x221(conv11out[221]),
.x222(conv11out[222]),
.x223(conv11out[223]),
.x224(conv11out[224]),
.x225(conv11out[225]),
.x226(conv11out[226]),
.x227(conv11out[227]),
.x228(conv11out[228]),
.x229(conv11out[229]),
.x230(conv11out[230]),
.x231(conv11out[231]),
.x232(conv11out[232]),
.x233(conv11out[233]),
.x234(conv11out[234]),
.x235(conv11out[235]),
.x236(conv11out[236]),
.x237(conv11out[237]),
.x238(conv11out[238]),
.x239(conv11out[239]),
.x240(conv11out[240]),
.x241(conv11out[241]),
.x242(conv11out[242]),
.x243(conv11out[243]),
.x244(conv11out[244]),
.x245(conv11out[245]),
.x246(conv11out[246]),
.x247(conv11out[247]),
.x248(conv11out[248]),
.x249(conv11out[249]),
.x250(conv11out[250]),
.x251(conv11out[251]),
.x252(conv11out[252]),
.x253(conv11out[253]),
.x254(conv11out[254]),
.x255(conv11out[255]),
.x256(conv11out[256]),
.x257(conv11out[257]),
.x258(conv11out[258]),
.x259(conv11out[259]),
.x260(conv11out[260]),
.x261(conv11out[261]),
.x262(conv11out[262]),
.x263(conv11out[263]),
.x264(conv11out[264]),
.x265(conv11out[265]),
.x266(conv11out[266]),
.x267(conv11out[267]),
.x268(conv11out[268]),
.x269(conv11out[269]),
.x270(conv11out[270]),
.x271(conv11out[271]),
.x272(conv11out[272]),
.x273(conv11out[273]),
.x274(conv11out[274]),
.x275(conv11out[275]),
.x276(conv11out[276]),
.x277(conv11out[277]),
.x278(conv11out[278]),
.x279(conv11out[279]),
.x280(conv11out[280]),
.x281(conv11out[281]),
.x282(conv11out[282]),
.x283(conv11out[283]),
.x284(conv11out[284]),
.x285(conv11out[285]),
.x286(conv11out[286]),
.x287(conv11out[287]),
.x288(conv11out[288]),
.x289(conv11out[289]),
.x290(conv11out[290]),
.x291(conv11out[291]),
.x292(conv11out[292]),
.x293(conv11out[293]),
.x294(conv11out[294]),
.x295(conv11out[295]),
.x296(conv11out[296]),
.x297(conv11out[297]),
.x298(conv11out[298]),
.x299(conv11out[299]),
.x300(conv11out[300]),
.x301(conv11out[301]),
.x302(conv11out[302]),
.x303(conv11out[303]),
.x304(conv11out[304]),
.x305(conv11out[305]),
.x306(conv11out[306]),
.x307(conv11out[307]),
.x308(conv11out[308]),
.x309(conv11out[309]),
.x310(conv11out[310]),
.x311(conv11out[311]),
.x312(conv11out[312]),
.x313(conv11out[313]),
.x314(conv11out[314]),
.x315(conv11out[315]),
.x316(conv11out[316]),
.x317(conv11out[317]),
.x318(conv11out[318]),
.x319(conv11out[319]),
.x320(conv11out[320]),
.x321(conv11out[321]),
.x322(conv11out[322]),
.x323(conv11out[323]),
.x324(conv11out[324]),
.x325(conv11out[325]),
.x326(conv11out[326]),
.x327(conv11out[327]),
.x328(conv11out[328]),
.x329(conv11out[329]),
.x330(conv11out[330]),
.x331(conv11out[331]),
.x332(conv11out[332]),
.x333(conv11out[333]),
.x334(conv11out[334]),
.x335(conv11out[335]),
.x336(conv11out[336]),
.x337(conv11out[337]),
.x338(conv11out[338]),
.x339(conv11out[339]),
.x340(conv11out[340]),
.x341(conv11out[341]),
.x342(conv11out[342]),
.x343(conv11out[343]),
.x344(conv11out[344]),
.x345(conv11out[345]),
.x346(conv11out[346]),
.x347(conv11out[347]),
.x348(conv11out[348]),
.x349(conv11out[349]),
.x350(conv11out[350]),
.x351(conv11out[351]),
.x352(conv11out[352]),
.x353(conv11out[353]),
.x354(conv11out[354]),
.x355(conv11out[355]),
.x356(conv11out[356]),
.x357(conv11out[357]),
.x358(conv11out[358]),
.x359(conv11out[359]),
.x360(conv11out[360]),
.x361(conv11out[361]),
.x362(conv11out[362]),
.x363(conv11out[363]),
.x364(conv11out[364]),
.x365(conv11out[365]),
.x366(conv11out[366]),
.x367(conv11out[367]),
.x368(conv11out[368]),
.x369(conv11out[369]),
.x370(conv11out[370]),
.x371(conv11out[371]),
.x372(conv11out[372]),
.x373(conv11out[373]),
.x374(conv11out[374]),
.x375(conv11out[375]),
.x376(conv11out[376]),
.x377(conv11out[377]),
.x378(conv11out[378]),
.x379(conv11out[379]),
.x380(conv11out[380]),
.x381(conv11out[381]),
.x382(conv11out[382]),
.x383(conv11out[383]),
.x384(conv11out[384]),
.x385(conv11out[385]),
.x386(conv11out[386]),
.x387(conv11out[387]),
.x388(conv11out[388]),
.x389(conv11out[389]),
.x390(conv11out[390]),
.x391(conv11out[391]),
.x392(conv11out[392]),
.x393(conv11out[393]),
.x394(conv11out[394]),
.x395(conv11out[395]),
.x396(conv11out[396]),
.x397(conv11out[397]),
.x398(conv11out[398]),
.x399(conv11out[399]),
.x400(conv11out[400]),
.x401(conv11out[401]),
.x402(conv11out[402]),
.x403(conv11out[403]),
.x404(conv11out[404]),
.x405(conv11out[405]),
.x406(conv11out[406]),
.x407(conv11out[407]),
.x408(conv11out[408]),
.x409(conv11out[409]),
.x410(conv11out[410]),
.x411(conv11out[411]),
.x412(conv11out[412]),
.x413(conv11out[413]),
.x414(conv11out[414]),
.x415(conv11out[415]),
.x416(conv11out[416]),
.x417(conv11out[417]),
.x418(conv11out[418]),
.x419(conv11out[419]),
.x420(conv11out[420]),
.x421(conv11out[421]),
.x422(conv11out[422]),
.x423(conv11out[423]),
.x424(conv11out[424]),
.x425(conv11out[425]),
.x426(conv11out[426]),
.x427(conv11out[427]),
.x428(conv11out[428]),
.x429(conv11out[429]),
.x430(conv11out[430]),
.x431(conv11out[431]),
.x432(conv11out[432]),
.x433(conv11out[433]),
.x434(conv11out[434]),
.x435(conv11out[435]),
.x436(conv11out[436]),
.x437(conv11out[437]),
.x438(conv11out[438]),
.x439(conv11out[439]),
.x440(conv11out[440]),
.x441(conv11out[441]),
.x442(conv11out[442]),
.x443(conv11out[443]),
.x444(conv11out[444]),
.x445(conv11out[445]),
.x446(conv11out[446]),
.x447(conv11out[447]),
.x448(conv11out[448]),
.x449(conv11out[449]),
.x450(conv11out[450]),
.x451(conv11out[451]),
.x452(conv11out[452]),
.x453(conv11out[453]),
.x454(conv11out[454]),
.x455(conv11out[455]),
.x456(conv11out[456]),
.x457(conv11out[457]),
.x458(conv11out[458]),
.x459(conv11out[459]),
.x460(conv11out[460]),
.x461(conv11out[461]),
.x462(conv11out[462]),
.x463(conv11out[463]),
.x464(conv11out[464]),
.x465(conv11out[465]),
.x466(conv11out[466]),
.x467(conv11out[467]),
.x468(conv11out[468]),
.x469(conv11out[469]),
.x470(conv11out[470]),
.x471(conv11out[471]),
.x472(conv11out[472]),
.x473(conv11out[473]),
.x474(conv11out[474]),
.x475(conv11out[475]),
.x476(conv11out[476]),
.x477(conv11out[477]),
.x478(conv11out[478]),
.x479(conv11out[479]),
.x480(conv11out[480]),
.x481(conv11out[481]),
.x482(conv11out[482]),
.x483(conv11out[483]),
.x484(conv11out[484]),
.x485(conv11out[485]),
.x486(conv11out[486]),
.x487(conv11out[487]),
.x488(conv11out[488]),
.x489(conv11out[489]),
.x490(conv11out[490]),
.x491(conv11out[491]),
.x492(conv11out[492]),
.x493(conv11out[493]),
.x494(conv11out[494]),
.x495(conv11out[495]),
.x496(conv11out[496]),
.x497(conv11out[497]),
.x498(conv11out[498]),
.x499(conv11out[499]),
.x500(conv11out[500]),
.x501(conv11out[501]),
.x502(conv11out[502]),
.x503(conv11out[503]),
.x504(conv11out[504]),
.x505(conv11out[505]),
.x506(conv11out[506]),
.x507(conv11out[507]),
.x508(conv11out[508]),
.x509(conv11out[509]),
.x510(conv11out[510]),
.x511(conv11out[511]),
.y0(conv21out[0]),
.y1(conv21out[1]),
.y2(conv21out[2]),
.y3(conv21out[3]),
.y4(conv21out[4]),
.y5(conv21out[5]),
.y6(conv21out[6]),
.y7(conv21out[7]),
.y8(conv21out[8]),
.y9(conv21out[9]),
.y10(conv21out[10]),
.y11(conv21out[11]),
.y12(conv21out[12]),
.y13(conv21out[13]),
.y14(conv21out[14]),
.y15(conv21out[15]),
.y16(conv21out[16]),
.y17(conv21out[17]),
.y18(conv21out[18]),
.y19(conv21out[19]),
.y20(conv21out[20]),
.y21(conv21out[21]),
.y22(conv21out[22]),
.y23(conv21out[23]),
.y24(conv21out[24]),
.y25(conv21out[25]),
.y26(conv21out[26]),
.y27(conv21out[27]),
.y28(conv21out[28]),
.y29(conv21out[29]),
.y30(conv21out[30]),
.y31(conv21out[31]),
.y32(conv21out[32]),
.y33(conv21out[33]),
.y34(conv21out[34]),
.y35(conv21out[35]),
.y36(conv21out[36]),
.y37(conv21out[37]),
.y38(conv21out[38]),
.y39(conv21out[39]),
.y40(conv21out[40]),
.y41(conv21out[41]),
.y42(conv21out[42]),
.y43(conv21out[43]),
.y44(conv21out[44]),
.y45(conv21out[45]),
.y46(conv21out[46]),
.y47(conv21out[47]),
.y48(conv21out[48]),
.y49(conv21out[49]),
.y50(conv21out[50]),
.y51(conv21out[51]),
.y52(conv21out[52]),
.y53(conv21out[53]),
.y54(conv21out[54]),
.y55(conv21out[55]),
.y56(conv21out[56]),
.y57(conv21out[57]),
.y58(conv21out[58]),
.y59(conv21out[59]),
.y60(conv21out[60]),
.y61(conv21out[61]),
.y62(conv21out[62]),
.y63(conv21out[63]),
.y64(conv21out[64]),
.y65(conv21out[65]),
.y66(conv21out[66]),
.y67(conv21out[67]),
.y68(conv21out[68]),
.y69(conv21out[69]),
.y70(conv21out[70]),
.y71(conv21out[71]),
.y72(conv21out[72]),
.y73(conv21out[73]),
.y74(conv21out[74]),
.y75(conv21out[75]),
.y76(conv21out[76]),
.y77(conv21out[77]),
.y78(conv21out[78]),
.y79(conv21out[79]),
.y80(conv21out[80]),
.y81(conv21out[81]),
.y82(conv21out[82]),
.y83(conv21out[83]),
.y84(conv21out[84]),
.y85(conv21out[85]),
.y86(conv21out[86]),
.y87(conv21out[87]),
.y88(conv21out[88]),
.y89(conv21out[89]),
.y90(conv21out[90]),
.y91(conv21out[91]),
.y92(conv21out[92]),
.y93(conv21out[93]),
.y94(conv21out[94]),
.y95(conv21out[95]),
.y96(conv21out[96]),
.y97(conv21out[97]),
.y98(conv21out[98]),
.y99(conv21out[99]),
.y100(conv21out[100]),
.y101(conv21out[101]),
.y102(conv21out[102]),
.y103(conv21out[103]),
.y104(conv21out[104]),
.y105(conv21out[105]),
.y106(conv21out[106]),
.y107(conv21out[107]),
.y108(conv21out[108]),
.y109(conv21out[109]),
.y110(conv21out[110]),
.y111(conv21out[111]),
.y112(conv21out[112]),
.y113(conv21out[113]),
.y114(conv21out[114]),
.y115(conv21out[115]),
.y116(conv21out[116]),
.y117(conv21out[117]),
.y118(conv21out[118]),
.y119(conv21out[119]),
.y120(conv21out[120]),
.y121(conv21out[121]),
.y122(conv21out[122]),
.y123(conv21out[123]),
.y124(conv21out[124]),
.y125(conv21out[125]),
.y126(conv21out[126]),
.y127(conv21out[127]),
.y128(conv21out[128]),
.y129(conv21out[129]),
.y130(conv21out[130]),
.y131(conv21out[131]),
.y132(conv21out[132]),
.y133(conv21out[133]),
.y134(conv21out[134]),
.y135(conv21out[135]),
.y136(conv21out[136]),
.y137(conv21out[137]),
.y138(conv21out[138]),
.y139(conv21out[139]),
.y140(conv21out[140]),
.y141(conv21out[141]),
.y142(conv21out[142]),
.y143(conv21out[143]),
.y144(conv21out[144]),
.y145(conv21out[145]),
.y146(conv21out[146]),
.y147(conv21out[147]),
.y148(conv21out[148]),
.y149(conv21out[149]),
.y150(conv21out[150]),
.y151(conv21out[151]),
.y152(conv21out[152]),
.y153(conv21out[153]),
.y154(conv21out[154]),
.y155(conv21out[155]),
.y156(conv21out[156]),
.y157(conv21out[157]),
.y158(conv21out[158]),
.y159(conv21out[159]),
.y160(conv21out[160]),
.y161(conv21out[161]),
.y162(conv21out[162]),
.y163(conv21out[163]),
.y164(conv21out[164]),
.y165(conv21out[165]),
.y166(conv21out[166]),
.y167(conv21out[167]),
.y168(conv21out[168]),
.y169(conv21out[169]),
.y170(conv21out[170]),
.y171(conv21out[171]),
.y172(conv21out[172]),
.y173(conv21out[173]),
.y174(conv21out[174]),
.y175(conv21out[175]),
.y176(conv21out[176]),
.y177(conv21out[177]),
.y178(conv21out[178]),
.y179(conv21out[179]),
.y180(conv21out[180]),
.y181(conv21out[181]),
.y182(conv21out[182]),
.y183(conv21out[183]),
.y184(conv21out[184]),
.y185(conv21out[185]),
.y186(conv21out[186]),
.y187(conv21out[187]),
.y188(conv21out[188]),
.y189(conv21out[189]),
.y190(conv21out[190]),
.y191(conv21out[191]),
.y192(conv21out[192]),
.y193(conv21out[193]),
.y194(conv21out[194]),
.y195(conv21out[195]),
.y196(conv21out[196]),
.y197(conv21out[197]),
.y198(conv21out[198]),
.y199(conv21out[199]),
.y200(conv21out[200]),
.y201(conv21out[201]),
.y202(conv21out[202]),
.y203(conv21out[203]),
.y204(conv21out[204]),
.y205(conv21out[205]),
.y206(conv21out[206]),
.y207(conv21out[207]),
.y208(conv21out[208]),
.y209(conv21out[209]),
.y210(conv21out[210]),
.y211(conv21out[211]),
.y212(conv21out[212]),
.y213(conv21out[213]),
.y214(conv21out[214]),
.y215(conv21out[215]),
.y216(conv21out[216]),
.y217(conv21out[217]),
.y218(conv21out[218]),
.y219(conv21out[219]),
.y220(conv21out[220]),
.y221(conv21out[221]),
.y222(conv21out[222]),
.y223(conv21out[223]),
.y224(conv21out[224]),
.y225(conv21out[225]),
.y226(conv21out[226]),
.y227(conv21out[227]),
.y228(conv21out[228]),
.y229(conv21out[229]),
.y230(conv21out[230]),
.y231(conv21out[231]),
.y232(conv21out[232]),
.y233(conv21out[233]),
.y234(conv21out[234]),
.y235(conv21out[235]),
.y236(conv21out[236]),
.y237(conv21out[237]),
.y238(conv21out[238]),
.y239(conv21out[239]),
.y240(conv21out[240]),
.y241(conv21out[241]),
.y242(conv21out[242]),
.y243(conv21out[243]),
.y244(conv21out[244]),
.y245(conv21out[245]),
.y246(conv21out[246]),
.y247(conv21out[247]),
.y248(conv21out[248]),
.y249(conv21out[249]),
.y250(conv21out[250]),
.y251(conv21out[251]),
.y252(conv21out[252]),
.y253(conv21out[253]),
.y254(conv21out[254]),
.y255(conv21out[255]),
.y256(conv21out[256]),
.y257(conv21out[257]),
.y258(conv21out[258]),
.y259(conv21out[259]),
.y260(conv21out[260]),
.y261(conv21out[261]),
.y262(conv21out[262]),
.y263(conv21out[263]),
.y264(conv21out[264]),
.y265(conv21out[265]),
.y266(conv21out[266]),
.y267(conv21out[267]),
.y268(conv21out[268]),
.y269(conv21out[269]),
.y270(conv21out[270]),
.y271(conv21out[271]),
.y272(conv21out[272]),
.y273(conv21out[273]),
.y274(conv21out[274]),
.y275(conv21out[275]),
.y276(conv21out[276]),
.y277(conv21out[277]),
.y278(conv21out[278]),
.y279(conv21out[279]),
.y280(conv21out[280]),
.y281(conv21out[281]),
.y282(conv21out[282]),
.y283(conv21out[283]),
.y284(conv21out[284]),
.y285(conv21out[285]),
.y286(conv21out[286]),
.y287(conv21out[287]) );
Conv22 conv22(.x0(conv11out[256]),
.x1(conv11out[257]),
.x2(conv11out[258]),
.x3(conv11out[259]),
.x4(conv11out[260]),
.x5(conv11out[261]),
.x6(conv11out[262]),
.x7(conv11out[263]),
.x8(conv11out[264]),
.x9(conv11out[265]),
.x10(conv11out[266]),
.x11(conv11out[267]),
.x12(conv11out[268]),
.x13(conv11out[269]),
.x14(conv11out[270]),
.x15(conv11out[271]),
.x16(conv11out[272]),
.x17(conv11out[273]),
.x18(conv11out[274]),
.x19(conv11out[275]),
.x20(conv11out[276]),
.x21(conv11out[277]),
.x22(conv11out[278]),
.x23(conv11out[279]),
.x24(conv11out[280]),
.x25(conv11out[281]),
.x26(conv11out[282]),
.x27(conv11out[283]),
.x28(conv11out[284]),
.x29(conv11out[285]),
.x30(conv11out[286]),
.x31(conv11out[287]),
.x32(conv11out[288]),
.x33(conv11out[289]),
.x34(conv11out[290]),
.x35(conv11out[291]),
.x36(conv11out[292]),
.x37(conv11out[293]),
.x38(conv11out[294]),
.x39(conv11out[295]),
.x40(conv11out[296]),
.x41(conv11out[297]),
.x42(conv11out[298]),
.x43(conv11out[299]),
.x44(conv11out[300]),
.x45(conv11out[301]),
.x46(conv11out[302]),
.x47(conv11out[303]),
.x48(conv11out[304]),
.x49(conv11out[305]),
.x50(conv11out[306]),
.x51(conv11out[307]),
.x52(conv11out[308]),
.x53(conv11out[309]),
.x54(conv11out[310]),
.x55(conv11out[311]),
.x56(conv11out[312]),
.x57(conv11out[313]),
.x58(conv11out[314]),
.x59(conv11out[315]),
.x60(conv11out[316]),
.x61(conv11out[317]),
.x62(conv11out[318]),
.x63(conv11out[319]),
.x64(conv11out[320]),
.x65(conv11out[321]),
.x66(conv11out[322]),
.x67(conv11out[323]),
.x68(conv11out[324]),
.x69(conv11out[325]),
.x70(conv11out[326]),
.x71(conv11out[327]),
.x72(conv11out[328]),
.x73(conv11out[329]),
.x74(conv11out[330]),
.x75(conv11out[331]),
.x76(conv11out[332]),
.x77(conv11out[333]),
.x78(conv11out[334]),
.x79(conv11out[335]),
.x80(conv11out[336]),
.x81(conv11out[337]),
.x82(conv11out[338]),
.x83(conv11out[339]),
.x84(conv11out[340]),
.x85(conv11out[341]),
.x86(conv11out[342]),
.x87(conv11out[343]),
.x88(conv11out[344]),
.x89(conv11out[345]),
.x90(conv11out[346]),
.x91(conv11out[347]),
.x92(conv11out[348]),
.x93(conv11out[349]),
.x94(conv11out[350]),
.x95(conv11out[351]),
.x96(conv11out[352]),
.x97(conv11out[353]),
.x98(conv11out[354]),
.x99(conv11out[355]),
.x100(conv11out[356]),
.x101(conv11out[357]),
.x102(conv11out[358]),
.x103(conv11out[359]),
.x104(conv11out[360]),
.x105(conv11out[361]),
.x106(conv11out[362]),
.x107(conv11out[363]),
.x108(conv11out[364]),
.x109(conv11out[365]),
.x110(conv11out[366]),
.x111(conv11out[367]),
.x112(conv11out[368]),
.x113(conv11out[369]),
.x114(conv11out[370]),
.x115(conv11out[371]),
.x116(conv11out[372]),
.x117(conv11out[373]),
.x118(conv11out[374]),
.x119(conv11out[375]),
.x120(conv11out[376]),
.x121(conv11out[377]),
.x122(conv11out[378]),
.x123(conv11out[379]),
.x124(conv11out[380]),
.x125(conv11out[381]),
.x126(conv11out[382]),
.x127(conv11out[383]),
.x128(conv11out[384]),
.x129(conv11out[385]),
.x130(conv11out[386]),
.x131(conv11out[387]),
.x132(conv11out[388]),
.x133(conv11out[389]),
.x134(conv11out[390]),
.x135(conv11out[391]),
.x136(conv11out[392]),
.x137(conv11out[393]),
.x138(conv11out[394]),
.x139(conv11out[395]),
.x140(conv11out[396]),
.x141(conv11out[397]),
.x142(conv11out[398]),
.x143(conv11out[399]),
.x144(conv11out[400]),
.x145(conv11out[401]),
.x146(conv11out[402]),
.x147(conv11out[403]),
.x148(conv11out[404]),
.x149(conv11out[405]),
.x150(conv11out[406]),
.x151(conv11out[407]),
.x152(conv11out[408]),
.x153(conv11out[409]),
.x154(conv11out[410]),
.x155(conv11out[411]),
.x156(conv11out[412]),
.x157(conv11out[413]),
.x158(conv11out[414]),
.x159(conv11out[415]),
.x160(conv11out[416]),
.x161(conv11out[417]),
.x162(conv11out[418]),
.x163(conv11out[419]),
.x164(conv11out[420]),
.x165(conv11out[421]),
.x166(conv11out[422]),
.x167(conv11out[423]),
.x168(conv11out[424]),
.x169(conv11out[425]),
.x170(conv11out[426]),
.x171(conv11out[427]),
.x172(conv11out[428]),
.x173(conv11out[429]),
.x174(conv11out[430]),
.x175(conv11out[431]),
.x176(conv11out[432]),
.x177(conv11out[433]),
.x178(conv11out[434]),
.x179(conv11out[435]),
.x180(conv11out[436]),
.x181(conv11out[437]),
.x182(conv11out[438]),
.x183(conv11out[439]),
.x184(conv11out[440]),
.x185(conv11out[441]),
.x186(conv11out[442]),
.x187(conv11out[443]),
.x188(conv11out[444]),
.x189(conv11out[445]),
.x190(conv11out[446]),
.x191(conv11out[447]),
.x192(conv11out[448]),
.x193(conv11out[449]),
.x194(conv11out[450]),
.x195(conv11out[451]),
.x196(conv11out[452]),
.x197(conv11out[453]),
.x198(conv11out[454]),
.x199(conv11out[455]),
.x200(conv11out[456]),
.x201(conv11out[457]),
.x202(conv11out[458]),
.x203(conv11out[459]),
.x204(conv11out[460]),
.x205(conv11out[461]),
.x206(conv11out[462]),
.x207(conv11out[463]),
.x208(conv11out[464]),
.x209(conv11out[465]),
.x210(conv11out[466]),
.x211(conv11out[467]),
.x212(conv11out[468]),
.x213(conv11out[469]),
.x214(conv11out[470]),
.x215(conv11out[471]),
.x216(conv11out[472]),
.x217(conv11out[473]),
.x218(conv11out[474]),
.x219(conv11out[475]),
.x220(conv11out[476]),
.x221(conv11out[477]),
.x222(conv11out[478]),
.x223(conv11out[479]),
.x224(conv11out[480]),
.x225(conv11out[481]),
.x226(conv11out[482]),
.x227(conv11out[483]),
.x228(conv11out[484]),
.x229(conv11out[485]),
.x230(conv11out[486]),
.x231(conv11out[487]),
.x232(conv11out[488]),
.x233(conv11out[489]),
.x234(conv11out[490]),
.x235(conv11out[491]),
.x236(conv11out[492]),
.x237(conv11out[493]),
.x238(conv11out[494]),
.x239(conv11out[495]),
.x240(conv11out[496]),
.x241(conv11out[497]),
.x242(conv11out[498]),
.x243(conv11out[499]),
.x244(conv11out[500]),
.x245(conv11out[501]),
.x246(conv11out[502]),
.x247(conv11out[503]),
.x248(conv11out[504]),
.x249(conv11out[505]),
.x250(conv11out[506]),
.x251(conv11out[507]),
.x252(conv11out[508]),
.x253(conv11out[509]),
.x254(conv11out[510]),
.x255(conv11out[511]),
.x256(conv11out[512]),
.x257(conv11out[513]),
.x258(conv11out[514]),
.x259(conv11out[515]),
.x260(conv11out[516]),
.x261(conv11out[517]),
.x262(conv11out[518]),
.x263(conv11out[519]),
.x264(conv11out[520]),
.x265(conv11out[521]),
.x266(conv11out[522]),
.x267(conv11out[523]),
.x268(conv11out[524]),
.x269(conv11out[525]),
.x270(conv11out[526]),
.x271(conv11out[527]),
.x272(conv11out[528]),
.x273(conv11out[529]),
.x274(conv11out[530]),
.x275(conv11out[531]),
.x276(conv11out[532]),
.x277(conv11out[533]),
.x278(conv11out[534]),
.x279(conv11out[535]),
.x280(conv11out[536]),
.x281(conv11out[537]),
.x282(conv11out[538]),
.x283(conv11out[539]),
.x284(conv11out[540]),
.x285(conv11out[541]),
.x286(conv11out[542]),
.x287(conv11out[543]),
.x288(conv11out[544]),
.x289(conv11out[545]),
.x290(conv11out[546]),
.x291(conv11out[547]),
.x292(conv11out[548]),
.x293(conv11out[549]),
.x294(conv11out[550]),
.x295(conv11out[551]),
.x296(conv11out[552]),
.x297(conv11out[553]),
.x298(conv11out[554]),
.x299(conv11out[555]),
.x300(conv11out[556]),
.x301(conv11out[557]),
.x302(conv11out[558]),
.x303(conv11out[559]),
.x304(conv11out[560]),
.x305(conv11out[561]),
.x306(conv11out[562]),
.x307(conv11out[563]),
.x308(conv11out[564]),
.x309(conv11out[565]),
.x310(conv11out[566]),
.x311(conv11out[567]),
.x312(conv11out[568]),
.x313(conv11out[569]),
.x314(conv11out[570]),
.x315(conv11out[571]),
.x316(conv11out[572]),
.x317(conv11out[573]),
.x318(conv11out[574]),
.x319(conv11out[575]),
.x320(conv11out[576]),
.x321(conv11out[577]),
.x322(conv11out[578]),
.x323(conv11out[579]),
.x324(conv11out[580]),
.x325(conv11out[581]),
.x326(conv11out[582]),
.x327(conv11out[583]),
.x328(conv11out[584]),
.x329(conv11out[585]),
.x330(conv11out[586]),
.x331(conv11out[587]),
.x332(conv11out[588]),
.x333(conv11out[589]),
.x334(conv11out[590]),
.x335(conv11out[591]),
.x336(conv11out[592]),
.x337(conv11out[593]),
.x338(conv11out[594]),
.x339(conv11out[595]),
.x340(conv11out[596]),
.x341(conv11out[597]),
.x342(conv11out[598]),
.x343(conv11out[599]),
.x344(conv11out[600]),
.x345(conv11out[601]),
.x346(conv11out[602]),
.x347(conv11out[603]),
.x348(conv11out[604]),
.x349(conv11out[605]),
.x350(conv11out[606]),
.x351(conv11out[607]),
.x352(conv11out[608]),
.x353(conv11out[609]),
.x354(conv11out[610]),
.x355(conv11out[611]),
.x356(conv11out[612]),
.x357(conv11out[613]),
.x358(conv11out[614]),
.x359(conv11out[615]),
.x360(conv11out[616]),
.x361(conv11out[617]),
.x362(conv11out[618]),
.x363(conv11out[619]),
.x364(conv11out[620]),
.x365(conv11out[621]),
.x366(conv11out[622]),
.x367(conv11out[623]),
.x368(conv11out[624]),
.x369(conv11out[625]),
.x370(conv11out[626]),
.x371(conv11out[627]),
.x372(conv11out[628]),
.x373(conv11out[629]),
.x374(conv11out[630]),
.x375(conv11out[631]),
.x376(conv11out[632]),
.x377(conv11out[633]),
.x378(conv11out[634]),
.x379(conv11out[635]),
.x380(conv11out[636]),
.x381(conv11out[637]),
.x382(conv11out[638]),
.x383(conv11out[639]),
.y0(conv22out[0]),
.y1(conv22out[1]),
.y2(conv22out[2]),
.y3(conv22out[3]),
.y4(conv22out[4]),
.y5(conv22out[5]),
.y6(conv22out[6]),
.y7(conv22out[7]),
.y8(conv22out[8]),
.y9(conv22out[9]),
.y10(conv22out[10]),
.y11(conv22out[11]),
.y12(conv22out[12]),
.y13(conv22out[13]),
.y14(conv22out[14]),
.y15(conv22out[15]),
.y16(conv22out[16]),
.y17(conv22out[17]),
.y18(conv22out[18]),
.y19(conv22out[19]),
.y20(conv22out[20]),
.y21(conv22out[21]),
.y22(conv22out[22]),
.y23(conv22out[23]),
.y24(conv22out[24]),
.y25(conv22out[25]),
.y26(conv22out[26]),
.y27(conv22out[27]),
.y28(conv22out[28]),
.y29(conv22out[29]),
.y30(conv22out[30]),
.y31(conv22out[31]),
.y32(conv22out[32]),
.y33(conv22out[33]),
.y34(conv22out[34]),
.y35(conv22out[35]),
.y36(conv22out[36]),
.y37(conv22out[37]),
.y38(conv22out[38]),
.y39(conv22out[39]),
.y40(conv22out[40]),
.y41(conv22out[41]),
.y42(conv22out[42]),
.y43(conv22out[43]),
.y44(conv22out[44]),
.y45(conv22out[45]),
.y46(conv22out[46]),
.y47(conv22out[47]),
.y48(conv22out[48]),
.y49(conv22out[49]),
.y50(conv22out[50]),
.y51(conv22out[51]),
.y52(conv22out[52]),
.y53(conv22out[53]),
.y54(conv22out[54]),
.y55(conv22out[55]),
.y56(conv22out[56]),
.y57(conv22out[57]),
.y58(conv22out[58]),
.y59(conv22out[59]),
.y60(conv22out[60]),
.y61(conv22out[61]),
.y62(conv22out[62]),
.y63(conv22out[63]),
.y64(conv22out[64]),
.y65(conv22out[65]),
.y66(conv22out[66]),
.y67(conv22out[67]),
.y68(conv22out[68]),
.y69(conv22out[69]),
.y70(conv22out[70]),
.y71(conv22out[71]),
.y72(conv22out[72]),
.y73(conv22out[73]),
.y74(conv22out[74]),
.y75(conv22out[75]),
.y76(conv22out[76]),
.y77(conv22out[77]),
.y78(conv22out[78]),
.y79(conv22out[79]),
.y80(conv22out[80]),
.y81(conv22out[81]),
.y82(conv22out[82]),
.y83(conv22out[83]),
.y84(conv22out[84]),
.y85(conv22out[85]),
.y86(conv22out[86]),
.y87(conv22out[87]),
.y88(conv22out[88]),
.y89(conv22out[89]),
.y90(conv22out[90]),
.y91(conv22out[91]),
.y92(conv22out[92]),
.y93(conv22out[93]),
.y94(conv22out[94]),
.y95(conv22out[95]),
.y96(conv22out[96]),
.y97(conv22out[97]),
.y98(conv22out[98]),
.y99(conv22out[99]),
.y100(conv22out[100]),
.y101(conv22out[101]),
.y102(conv22out[102]),
.y103(conv22out[103]),
.y104(conv22out[104]),
.y105(conv22out[105]),
.y106(conv22out[106]),
.y107(conv22out[107]),
.y108(conv22out[108]),
.y109(conv22out[109]),
.y110(conv22out[110]),
.y111(conv22out[111]),
.y112(conv22out[112]),
.y113(conv22out[113]),
.y114(conv22out[114]),
.y115(conv22out[115]),
.y116(conv22out[116]),
.y117(conv22out[117]),
.y118(conv22out[118]),
.y119(conv22out[119]),
.y120(conv22out[120]),
.y121(conv22out[121]),
.y122(conv22out[122]),
.y123(conv22out[123]),
.y124(conv22out[124]),
.y125(conv22out[125]),
.y126(conv22out[126]),
.y127(conv22out[127]),
.y128(conv22out[128]),
.y129(conv22out[129]),
.y130(conv22out[130]),
.y131(conv22out[131]),
.y132(conv22out[132]),
.y133(conv22out[133]),
.y134(conv22out[134]),
.y135(conv22out[135]),
.y136(conv22out[136]),
.y137(conv22out[137]),
.y138(conv22out[138]),
.y139(conv22out[139]),
.y140(conv22out[140]),
.y141(conv22out[141]),
.y142(conv22out[142]),
.y143(conv22out[143]),
.y144(conv22out[144]),
.y145(conv22out[145]),
.y146(conv22out[146]),
.y147(conv22out[147]),
.y148(conv22out[148]),
.y149(conv22out[149]),
.y150(conv22out[150]),
.y151(conv22out[151]),
.y152(conv22out[152]),
.y153(conv22out[153]),
.y154(conv22out[154]),
.y155(conv22out[155]),
.y156(conv22out[156]),
.y157(conv22out[157]),
.y158(conv22out[158]),
.y159(conv22out[159]),
.y160(conv22out[160]),
.y161(conv22out[161]),
.y162(conv22out[162]),
.y163(conv22out[163]),
.y164(conv22out[164]),
.y165(conv22out[165]),
.y166(conv22out[166]),
.y167(conv22out[167]),
.y168(conv22out[168]),
.y169(conv22out[169]),
.y170(conv22out[170]),
.y171(conv22out[171]),
.y172(conv22out[172]),
.y173(conv22out[173]),
.y174(conv22out[174]),
.y175(conv22out[175]),
.y176(conv22out[176]),
.y177(conv22out[177]),
.y178(conv22out[178]),
.y179(conv22out[179]),
.y180(conv22out[180]),
.y181(conv22out[181]),
.y182(conv22out[182]),
.y183(conv22out[183]),
.y184(conv22out[184]),
.y185(conv22out[185]),
.y186(conv22out[186]),
.y187(conv22out[187]),
.y188(conv22out[188]),
.y189(conv22out[189]),
.y190(conv22out[190]),
.y191(conv22out[191]),
.y192(conv22out[192]),
.y193(conv22out[193]),
.y194(conv22out[194]),
.y195(conv22out[195]),
.y196(conv22out[196]),
.y197(conv22out[197]),
.y198(conv22out[198]),
.y199(conv22out[199]),
.y200(conv22out[200]),
.y201(conv22out[201]),
.y202(conv22out[202]),
.y203(conv22out[203]),
.y204(conv22out[204]),
.y205(conv22out[205]),
.y206(conv22out[206]),
.y207(conv22out[207]) );
Dense1 dense1(.x0(conv21out[0]),
.x1(conv21out[1]),
.x2(conv21out[2]),
.x3(conv21out[3]),
.x4(conv21out[4]),
.x5(conv21out[5]),
.x6(conv21out[6]),
.x7(conv21out[7]),
.x8(conv21out[8]),
.x9(conv21out[9]),
.x10(conv21out[10]),
.x11(conv21out[11]),
.x12(conv21out[12]),
.x13(conv21out[13]),
.x14(conv21out[14]),
.x15(conv21out[15]),
.x16(conv21out[16]),
.x17(conv21out[17]),
.x18(conv21out[18]),
.x19(conv21out[19]),
.x20(conv21out[20]),
.x21(conv21out[21]),
.x22(conv21out[22]),
.x23(conv21out[23]),
.x24(conv21out[24]),
.x25(conv21out[25]),
.x26(conv21out[26]),
.x27(conv21out[27]),
.x28(conv21out[28]),
.x29(conv21out[29]),
.x30(conv21out[30]),
.x31(conv21out[31]),
.x32(conv21out[32]),
.x33(conv21out[33]),
.x34(conv21out[34]),
.x35(conv21out[35]),
.x36(conv21out[36]),
.x37(conv21out[37]),
.x38(conv21out[38]),
.x39(conv21out[39]),
.x40(conv21out[40]),
.x41(conv21out[41]),
.x42(conv21out[42]),
.x43(conv21out[43]),
.x44(conv21out[44]),
.x45(conv21out[45]),
.x46(conv21out[46]),
.x47(conv21out[47]),
.x48(conv21out[48]),
.x49(conv21out[49]),
.x50(conv21out[50]),
.x51(conv21out[51]),
.x52(conv21out[52]),
.x53(conv21out[53]),
.x54(conv21out[54]),
.x55(conv21out[55]),
.x56(conv21out[56]),
.x57(conv21out[57]),
.x58(conv21out[58]),
.x59(conv21out[59]),
.x60(conv21out[60]),
.x61(conv21out[61]),
.x62(conv21out[62]),
.x63(conv21out[63]),
.x64(conv21out[64]),
.x65(conv21out[65]),
.x66(conv21out[66]),
.x67(conv21out[67]),
.x68(conv21out[68]),
.x69(conv21out[69]),
.x70(conv21out[70]),
.x71(conv21out[71]),
.x72(conv21out[72]),
.x73(conv21out[73]),
.x74(conv21out[74]),
.x75(conv21out[75]),
.x76(conv21out[76]),
.x77(conv21out[77]),
.x78(conv21out[78]),
.x79(conv21out[79]),
.x80(conv21out[80]),
.x81(conv21out[81]),
.x82(conv21out[82]),
.x83(conv21out[83]),
.x84(conv21out[84]),
.x85(conv21out[85]),
.x86(conv21out[86]),
.x87(conv21out[87]),
.x88(conv21out[88]),
.x89(conv21out[89]),
.x90(conv21out[90]),
.x91(conv21out[91]),
.x92(conv21out[92]),
.x93(conv21out[93]),
.x94(conv21out[94]),
.x95(conv21out[95]),
.x96(conv21out[96]),
.x97(conv21out[97]),
.x98(conv21out[98]),
.x99(conv21out[99]),
.x100(conv21out[100]),
.x101(conv21out[101]),
.x102(conv21out[102]),
.x103(conv21out[103]),
.x104(conv21out[104]),
.x105(conv21out[105]),
.x106(conv21out[106]),
.x107(conv21out[107]),
.x108(conv21out[108]),
.x109(conv21out[109]),
.x110(conv21out[110]),
.x111(conv21out[111]),
.x112(conv21out[112]),
.x113(conv21out[113]),
.x114(conv21out[114]),
.x115(conv21out[115]),
.x116(conv21out[116]),
.x117(conv21out[117]),
.x118(conv21out[118]),
.x119(conv21out[119]),
.x120(conv21out[120]),
.x121(conv21out[121]),
.x122(conv21out[122]),
.x123(conv21out[123]),
.x124(conv21out[124]),
.x125(conv21out[125]),
.x126(conv21out[126]),
.x127(conv21out[127]),
.x128(conv21out[128]),
.x129(conv21out[129]),
.x130(conv21out[130]),
.x131(conv21out[131]),
.x132(conv21out[132]),
.x133(conv21out[133]),
.x134(conv21out[134]),
.x135(conv21out[135]),
.x136(conv21out[136]),
.x137(conv21out[137]),
.x138(conv21out[138]),
.x139(conv21out[139]),
.x140(conv21out[140]),
.x141(conv21out[141]),
.x142(conv21out[142]),
.x143(conv21out[143]),
.x144(conv21out[144]),
.x145(conv21out[145]),
.x146(conv21out[146]),
.x147(conv21out[147]),
.x148(conv21out[148]),
.x149(conv21out[149]),
.x150(conv21out[150]),
.x151(conv21out[151]),
.x152(conv21out[152]),
.x153(conv21out[153]),
.x154(conv21out[154]),
.x155(conv21out[155]),
.x156(conv21out[156]),
.x157(conv21out[157]),
.x158(conv21out[158]),
.x159(conv21out[159]),
.x160(conv21out[160]),
.x161(conv21out[161]),
.x162(conv21out[162]),
.x163(conv21out[163]),
.x164(conv21out[164]),
.x165(conv21out[165]),
.x166(conv21out[166]),
.x167(conv21out[167]),
.x168(conv21out[168]),
.x169(conv21out[169]),
.x170(conv21out[170]),
.x171(conv21out[171]),
.x172(conv21out[172]),
.x173(conv21out[173]),
.x174(conv21out[174]),
.x175(conv21out[175]),
.x176(conv21out[176]),
.x177(conv21out[177]),
.x178(conv21out[178]),
.x179(conv21out[179]),
.x180(conv21out[180]),
.x181(conv21out[181]),
.x182(conv21out[182]),
.x183(conv21out[183]),
.x184(conv21out[184]),
.x185(conv21out[185]),
.x186(conv21out[186]),
.x187(conv21out[187]),
.x188(conv21out[188]),
.x189(conv21out[189]),
.x190(conv21out[190]),
.x191(conv21out[191]),
.x192(conv21out[192]),
.x193(conv21out[193]),
.x194(conv21out[194]),
.x195(conv21out[195]),
.x196(conv21out[196]),
.x197(conv21out[197]),
.x198(conv21out[198]),
.x199(conv21out[199]),
.x200(conv21out[200]),
.x201(conv21out[201]),
.x202(conv21out[202]),
.x203(conv21out[203]),
.x204(conv21out[204]),
.x205(conv21out[205]),
.x206(conv21out[206]),
.x207(conv21out[207]),
.x208(conv21out[208]),
.x209(conv21out[209]),
.x210(conv21out[210]),
.x211(conv21out[211]),
.x212(conv21out[212]),
.x213(conv21out[213]),
.x214(conv21out[214]),
.x215(conv21out[215]),
.x216(conv21out[216]),
.x217(conv21out[217]),
.x218(conv21out[218]),
.x219(conv21out[219]),
.x220(conv21out[220]),
.x221(conv21out[221]),
.x222(conv21out[222]),
.x223(conv21out[223]),
.x224(conv21out[224]),
.x225(conv21out[225]),
.x226(conv21out[226]),
.x227(conv21out[227]),
.x228(conv21out[228]),
.x229(conv21out[229]),
.x230(conv21out[230]),
.x231(conv21out[231]),
.x232(conv21out[232]),
.x233(conv21out[233]),
.x234(conv21out[234]),
.x235(conv21out[235]),
.x236(conv21out[236]),
.x237(conv21out[237]),
.x238(conv21out[238]),
.x239(conv21out[239]),
.x240(conv21out[240]),
.x241(conv21out[241]),
.x242(conv21out[242]),
.x243(conv21out[243]),
.x244(conv21out[244]),
.x245(conv21out[245]),
.x246(conv21out[246]),
.x247(conv21out[247]),
.x248(conv21out[248]),
.x249(conv21out[249]),
.x250(conv21out[250]),
.x251(conv21out[251]),
.x252(conv21out[252]),
.x253(conv21out[253]),
.x254(conv21out[254]),
.x255(conv21out[255]),
.x256(conv21out[256]),
.x257(conv21out[257]),
.x258(conv21out[258]),
.x259(conv21out[259]),
.x260(conv21out[260]),
.x261(conv21out[261]),
.x262(conv21out[262]),
.x263(conv21out[263]),
.x264(conv21out[264]),
.x265(conv21out[265]),
.x266(conv21out[266]),
.x267(conv21out[267]),
.x268(conv21out[268]),
.x269(conv21out[269]),
.x270(conv21out[270]),
.x271(conv21out[271]),
.x272(conv21out[272]),
.x273(conv21out[273]),
.x274(conv21out[274]),
.x275(conv21out[275]),
.x276(conv21out[276]),
.x277(conv21out[277]),
.x278(conv21out[278]),
.x279(conv21out[279]),
.x280(conv21out[280]),
.x281(conv21out[281]),
.x282(conv21out[282]),
.x283(conv21out[283]),
.x284(conv21out[284]),
.x285(conv21out[285]),
.x286(conv21out[286]),
.x287(conv21out[287]),
.x288(conv22out[0]),
.x289(conv22out[1]),
.x290(conv22out[2]),
.x291(conv22out[3]),
.x292(conv22out[4]),
.x293(conv22out[5]),
.x294(conv22out[6]),
.x295(conv22out[7]),
.x296(conv22out[8]),
.x297(conv22out[9]),
.x298(conv22out[10]),
.x299(conv22out[11]),
.x300(conv22out[12]),
.x301(conv22out[13]),
.x302(conv22out[14]),
.x303(conv22out[15]),
.x304(conv22out[16]),
.x305(conv22out[17]),
.x306(conv22out[18]),
.x307(conv22out[19]),
.x308(conv22out[20]),
.x309(conv22out[21]),
.x310(conv22out[22]),
.x311(conv22out[23]),
.x312(conv22out[24]),
.x313(conv22out[25]),
.x314(conv22out[26]),
.x315(conv22out[27]),
.x316(conv22out[28]),
.x317(conv22out[29]),
.x318(conv22out[30]),
.x319(conv22out[31]),
.x320(conv22out[32]),
.x321(conv22out[33]),
.x322(conv22out[34]),
.x323(conv22out[35]),
.x324(conv22out[36]),
.x325(conv22out[37]),
.x326(conv22out[38]),
.x327(conv22out[39]),
.x328(conv22out[40]),
.x329(conv22out[41]),
.x330(conv22out[42]),
.x331(conv22out[43]),
.x332(conv22out[44]),
.x333(conv22out[45]),
.x334(conv22out[46]),
.x335(conv22out[47]),
.x336(conv22out[48]),
.x337(conv22out[49]),
.x338(conv22out[50]),
.x339(conv22out[51]),
.x340(conv22out[52]),
.x341(conv22out[53]),
.x342(conv22out[54]),
.x343(conv22out[55]),
.x344(conv22out[56]),
.x345(conv22out[57]),
.x346(conv22out[58]),
.x347(conv22out[59]),
.x348(conv22out[60]),
.x349(conv22out[61]),
.x350(conv22out[62]),
.x351(conv22out[63]),
.x352(conv22out[64]),
.x353(conv22out[65]),
.x354(conv22out[66]),
.x355(conv22out[67]),
.x356(conv22out[68]),
.x357(conv22out[69]),
.x358(conv22out[70]),
.x359(conv22out[71]),
.x360(conv22out[72]),
.x361(conv22out[73]),
.x362(conv22out[74]),
.x363(conv22out[75]),
.x364(conv22out[76]),
.x365(conv22out[77]),
.x366(conv22out[78]),
.x367(conv22out[79]),
.x368(conv22out[80]),
.x369(conv22out[81]),
.x370(conv22out[82]),
.x371(conv22out[83]),
.x372(conv22out[84]),
.x373(conv22out[85]),
.x374(conv22out[86]),
.x375(conv22out[87]),
.x376(conv22out[88]),
.x377(conv22out[89]),
.x378(conv22out[90]),
.x379(conv22out[91]),
.x380(conv22out[92]),
.x381(conv22out[93]),
.x382(conv22out[94]),
.x383(conv22out[95]),
.x384(conv22out[96]),
.x385(conv22out[97]),
.x386(conv22out[98]),
.x387(conv22out[99]),
.x388(conv22out[100]),
.x389(conv22out[101]),
.x390(conv22out[102]),
.x391(conv22out[103]),
.x392(conv22out[104]),
.x393(conv22out[105]),
.x394(conv22out[106]),
.x395(conv22out[107]),
.x396(conv22out[108]),
.x397(conv22out[109]),
.x398(conv22out[110]),
.x399(conv22out[111]),
.x400(conv22out[112]),
.x401(conv22out[113]),
.x402(conv22out[114]),
.x403(conv22out[115]),
.x404(conv22out[116]),
.x405(conv22out[117]),
.x406(conv22out[118]),
.x407(conv22out[119]),
.x408(conv22out[120]),
.x409(conv22out[121]),
.x410(conv22out[122]),
.x411(conv22out[123]),
.x412(conv22out[124]),
.x413(conv22out[125]),
.x414(conv22out[126]),
.x415(conv22out[127]),
.x416(conv22out[128]),
.x417(conv22out[129]),
.x418(conv22out[130]),
.x419(conv22out[131]),
.x420(conv22out[132]),
.x421(conv22out[133]),
.x422(conv22out[134]),
.x423(conv22out[135]),
.x424(conv22out[136]),
.x425(conv22out[137]),
.x426(conv22out[138]),
.x427(conv22out[139]),
.x428(conv22out[140]),
.x429(conv22out[141]),
.x430(conv22out[142]),
.x431(conv22out[143]),
.x432(conv22out[144]),
.x433(conv22out[145]),
.x434(conv22out[146]),
.x435(conv22out[147]),
.x436(conv22out[148]),
.x437(conv22out[149]),
.x438(conv22out[150]),
.x439(conv22out[151]),
.x440(conv22out[152]),
.x441(conv22out[153]),
.x442(conv22out[154]),
.x443(conv22out[155]),
.x444(conv22out[156]),
.x445(conv22out[157]),
.x446(conv22out[158]),
.x447(conv22out[159]),
.x448(conv22out[160]),
.x449(conv22out[161]),
.x450(conv22out[162]),
.x451(conv22out[163]),
.x452(conv22out[164]),
.x453(conv22out[165]),
.x454(conv22out[166]),
.x455(conv22out[167]),
.x456(conv22out[168]),
.x457(conv22out[169]),
.x458(conv22out[170]),
.x459(conv22out[171]),
.x460(conv22out[172]),
.x461(conv22out[173]),
.x462(conv22out[174]),
.x463(conv22out[175]),
.x464(conv22out[176]),
.x465(conv22out[177]),
.x466(conv22out[178]),
.x467(conv22out[179]),
.x468(conv22out[180]),
.x469(conv22out[181]),
.x470(conv22out[182]),
.x471(conv22out[183]),
.x472(conv22out[184]),
.x473(conv22out[185]),
.x474(conv22out[186]),
.x475(conv22out[187]),
.x476(conv22out[188]),
.x477(conv22out[189]),
.x478(conv22out[190]),
.x479(conv22out[191]),
.x480(conv22out[192]),
.x481(conv22out[193]),
.x482(conv22out[194]),
.x483(conv22out[195]),
.x484(conv22out[196]),
.x485(conv22out[197]),
.x486(conv22out[198]),
.x487(conv22out[199]),
.x488(conv22out[200]),
.x489(conv22out[201]),
.x490(conv22out[202]),
.x491(conv22out[203]),
.x492(conv22out[204]),
.x493(conv22out[205]),
.x494(conv22out[206]),
.x495(conv22out[207]),
.y0(dense1out[0]),
.y1(dense1out[1]),
.y2(dense1out[2]),
.y3(dense1out[3]),
.y4(dense1out[4]),
.y5(dense1out[5]),
.y6(dense1out[6]),
.y7(dense1out[7]),
.y8(dense1out[8]),
.y9(dense1out[9]),
.y10(dense1out[10]),
.y11(dense1out[11]),
.y12(dense1out[12]),
.y13(dense1out[13]),
.y14(dense1out[14]),
.y15(dense1out[15]),
.y16(dense1out[16]),
.y17(dense1out[17]),
.y18(dense1out[18]),
.y19(dense1out[19]) );
Dense dense(.x0(dense1out[0]),
.x1(dense1out[1]),
.x2(dense1out[2]),
.x3(dense1out[3]),
.x4(dense1out[4]),
.x5(dense1out[5]),
.x6(dense1out[6]),
.x7(dense1out[7]),
.x8(dense1out[8]),
.x9(dense1out[9]),
.x10(dense1out[10]),
.x11(dense1out[11]),
.x12(dense1out[12]),
.x13(dense1out[13]),
.x14(dense1out[14]),
.x15(dense1out[15]),
.x16(dense1out[16]),
.x17(dense1out[17]),
.x18(dense1out[18]),
.x19(dense1out[19]),
.y(y));
endmodule