module Dense1(
input [4:0] x0 ,
input [4:0] x1 ,
input [4:0] x2 ,
input [4:0] x3 ,
input [4:0] x4 ,
input [4:0] x5 ,
input [4:0] x6 ,
input [4:0] x7 ,
input [4:0] x8 ,
input [4:0] x9 ,
input [4:0] x10 ,
input [4:0] x11 ,
input [4:0] x12 ,
input [4:0] x13 ,
input [4:0] x14 ,
input [4:0] x15 ,
input [4:0] x16 ,
input [4:0] x17 ,
input [4:0] x18 ,
input [4:0] x19 ,
input [4:0] x20 ,
input [4:0] x21 ,
input [4:0] x22 ,
input [4:0] x23 ,
input [4:0] x24 ,
input [4:0] x25 ,
input [4:0] x26 ,
input [4:0] x27 ,
input [4:0] x28 ,
input [4:0] x29 ,
input [4:0] x30 ,
input [4:0] x31 ,
input [4:0] x32 ,
input [4:0] x33 ,
input [4:0] x34 ,
input [4:0] x35 ,
input [4:0] x36 ,
input [4:0] x37 ,
input [4:0] x38 ,
input [4:0] x39 ,
input [4:0] x40 ,
input [4:0] x41 ,
input [4:0] x42 ,
input [4:0] x43 ,
input [4:0] x44 ,
input [4:0] x45 ,
input [4:0] x46 ,
input [4:0] x47 ,
input [4:0] x48 ,
input [4:0] x49 ,
input [4:0] x50 ,
input [4:0] x51 ,
input [4:0] x52 ,
input [4:0] x53 ,
input [4:0] x54 ,
input [4:0] x55 ,
input [4:0] x56 ,
input [4:0] x57 ,
input [4:0] x58 ,
input [4:0] x59 ,
input [4:0] x60 ,
input [4:0] x61 ,
input [4:0] x62 ,
input [4:0] x63 ,
input [4:0] x64 ,
input [4:0] x65 ,
input [4:0] x66 ,
input [4:0] x67 ,
input [4:0] x68 ,
input [4:0] x69 ,
input [4:0] x70 ,
input [4:0] x71 ,
input [4:0] x72 ,
input [4:0] x73 ,
input [4:0] x74 ,
input [4:0] x75 ,
input [4:0] x76 ,
input [4:0] x77 ,
input [4:0] x78 ,
input [4:0] x79 ,
input [4:0] x80 ,
input [4:0] x81 ,
input [4:0] x82 ,
input [4:0] x83 ,
input [4:0] x84 ,
input [4:0] x85 ,
input [4:0] x86 ,
input [4:0] x87 ,
input [4:0] x88 ,
input [4:0] x89 ,
input [4:0] x90 ,
input [4:0] x91 ,
input [4:0] x92 ,
input [4:0] x93 ,
input [4:0] x94 ,
input [4:0] x95 ,
input [4:0] x96 ,
input [4:0] x97 ,
input [4:0] x98 ,
input [4:0] x99 ,
input [4:0] x100 ,
input [4:0] x101 ,
input [4:0] x102 ,
input [4:0] x103 ,
input [4:0] x104 ,
input [4:0] x105 ,
input [4:0] x106 ,
input [4:0] x107 ,
input [4:0] x108 ,
input [4:0] x109 ,
input [4:0] x110 ,
input [4:0] x111 ,
input [4:0] x112 ,
input [4:0] x113 ,
input [4:0] x114 ,
input [4:0] x115 ,
input [4:0] x116 ,
input [4:0] x117 ,
input [4:0] x118 ,
input [4:0] x119 ,
input [4:0] x120 ,
input [4:0] x121 ,
input [4:0] x122 ,
input [4:0] x123 ,
input [4:0] x124 ,
input [4:0] x125 ,
input [4:0] x126 ,
input [4:0] x127 ,
input [4:0] x128 ,
input [4:0] x129 ,
input [4:0] x130 ,
input [4:0] x131 ,
input [4:0] x132 ,
input [4:0] x133 ,
input [4:0] x134 ,
input [4:0] x135 ,
input [4:0] x136 ,
input [4:0] x137 ,
input [4:0] x138 ,
input [4:0] x139 ,
input [4:0] x140 ,
input [4:0] x141 ,
input [4:0] x142 ,
input [4:0] x143 ,
input [4:0] x144 ,
input [4:0] x145 ,
input [4:0] x146 ,
input [4:0] x147 ,
input [4:0] x148 ,
input [4:0] x149 ,
input [4:0] x150 ,
input [4:0] x151 ,
input [4:0] x152 ,
input [4:0] x153 ,
input [4:0] x154 ,
input [4:0] x155 ,
input [4:0] x156 ,
input [4:0] x157 ,
input [4:0] x158 ,
input [4:0] x159 ,
input [4:0] x160 ,
input [4:0] x161 ,
input [4:0] x162 ,
input [4:0] x163 ,
input [4:0] x164 ,
input [4:0] x165 ,
input [4:0] x166 ,
input [4:0] x167 ,
input [4:0] x168 ,
input [4:0] x169 ,
input [4:0] x170 ,
input [4:0] x171 ,
input [4:0] x172 ,
input [4:0] x173 ,
input [4:0] x174 ,
input [4:0] x175 ,
input [4:0] x176 ,
input [4:0] x177 ,
input [4:0] x178 ,
input [4:0] x179 ,
input [4:0] x180 ,
input [4:0] x181 ,
input [4:0] x182 ,
input [4:0] x183 ,
input [4:0] x184 ,
input [4:0] x185 ,
input [4:0] x186 ,
input [4:0] x187 ,
input [4:0] x188 ,
input [4:0] x189 ,
input [4:0] x190 ,
input [4:0] x191 ,
input [4:0] x192 ,
input [4:0] x193 ,
input [4:0] x194 ,
input [4:0] x195 ,
input [4:0] x196 ,
input [4:0] x197 ,
input [4:0] x198 ,
input [4:0] x199 ,
input [4:0] x200 ,
input [4:0] x201 ,
input [4:0] x202 ,
input [4:0] x203 ,
input [4:0] x204 ,
input [4:0] x205 ,
input [4:0] x206 ,
input [4:0] x207 ,
input [4:0] x208 ,
input [4:0] x209 ,
input [4:0] x210 ,
input [4:0] x211 ,
input [4:0] x212 ,
input [4:0] x213 ,
input [4:0] x214 ,
input [4:0] x215 ,
input [4:0] x216 ,
input [4:0] x217 ,
input [4:0] x218 ,
input [4:0] x219 ,
input [4:0] x220 ,
input [4:0] x221 ,
input [4:0] x222 ,
input [4:0] x223 ,
input [4:0] x224 ,
input [4:0] x225 ,
input [4:0] x226 ,
input [4:0] x227 ,
input [4:0] x228 ,
input [4:0] x229 ,
input [4:0] x230 ,
input [4:0] x231 ,
input [4:0] x232 ,
input [4:0] x233 ,
input [4:0] x234 ,
input [4:0] x235 ,
input [4:0] x236 ,
input [4:0] x237 ,
input [4:0] x238 ,
input [4:0] x239 ,
input [4:0] x240 ,
input [4:0] x241 ,
input [4:0] x242 ,
input [4:0] x243 ,
input [4:0] x244 ,
input [4:0] x245 ,
input [4:0] x246 ,
input [4:0] x247 ,
input [4:0] x248 ,
input [4:0] x249 ,
input [4:0] x250 ,
input [4:0] x251 ,
input [4:0] x252 ,
input [4:0] x253 ,
input [4:0] x254 ,
input [4:0] x255 ,
input [4:0] x256 ,
input [4:0] x257 ,
input [4:0] x258 ,
input [4:0] x259 ,
input [4:0] x260 ,
input [4:0] x261 ,
input [4:0] x262 ,
input [4:0] x263 ,
input [4:0] x264 ,
input [4:0] x265 ,
input [4:0] x266 ,
input [4:0] x267 ,
input [4:0] x268 ,
input [4:0] x269 ,
input [4:0] x270 ,
input [4:0] x271 ,
input [4:0] x272 ,
input [4:0] x273 ,
input [4:0] x274 ,
input [4:0] x275 ,
input [4:0] x276 ,
input [4:0] x277 ,
input [4:0] x278 ,
input [4:0] x279 ,
input [4:0] x280 ,
input [4:0] x281 ,
input [4:0] x282 ,
input [4:0] x283 ,
input [4:0] x284 ,
input [4:0] x285 ,
input [4:0] x286 ,
input [4:0] x287 ,
input [4:0] x288 ,
input [4:0] x289 ,
input [4:0] x290 ,
input [4:0] x291 ,
input [4:0] x292 ,
input [4:0] x293 ,
input [4:0] x294 ,
input [4:0] x295 ,
input [4:0] x296 ,
input [4:0] x297 ,
input [4:0] x298 ,
input [4:0] x299 ,
input [4:0] x300 ,
input [4:0] x301 ,
input [4:0] x302 ,
input [4:0] x303 ,
input [4:0] x304 ,
input [4:0] x305 ,
input [4:0] x306 ,
input [4:0] x307 ,
input [4:0] x308 ,
input [4:0] x309 ,
input [4:0] x310 ,
input [4:0] x311 ,
input [4:0] x312 ,
input [4:0] x313 ,
input [4:0] x314 ,
input [4:0] x315 ,
input [4:0] x316 ,
input [4:0] x317 ,
input [4:0] x318 ,
input [4:0] x319 ,
input [4:0] x320 ,
input [4:0] x321 ,
input [4:0] x322 ,
input [4:0] x323 ,
input [4:0] x324 ,
input [4:0] x325 ,
input [4:0] x326 ,
input [4:0] x327 ,
input [4:0] x328 ,
input [4:0] x329 ,
input [4:0] x330 ,
input [4:0] x331 ,
input [4:0] x332 ,
input [4:0] x333 ,
input [4:0] x334 ,
input [4:0] x335 ,
input [4:0] x336 ,
input [4:0] x337 ,
input [4:0] x338 ,
input [4:0] x339 ,
input [4:0] x340 ,
input [4:0] x341 ,
input [4:0] x342 ,
input [4:0] x343 ,
input [4:0] x344 ,
input [4:0] x345 ,
input [4:0] x346 ,
input [4:0] x347 ,
input [4:0] x348 ,
input [4:0] x349 ,
input [4:0] x350 ,
input [4:0] x351 ,
input [4:0] x352 ,
input [4:0] x353 ,
input [4:0] x354 ,
input [4:0] x355 ,
input [4:0] x356 ,
input [4:0] x357 ,
input [4:0] x358 ,
input [4:0] x359 ,
input [4:0] x360 ,
input [4:0] x361 ,
input [4:0] x362 ,
input [4:0] x363 ,
input [4:0] x364 ,
input [4:0] x365 ,
input [4:0] x366 ,
input [4:0] x367 ,
input [4:0] x368 ,
input [4:0] x369 ,
input [4:0] x370 ,
input [4:0] x371 ,
input [4:0] x372 ,
input [4:0] x373 ,
input [4:0] x374 ,
input [4:0] x375 ,
input [4:0] x376 ,
input [4:0] x377 ,
input [4:0] x378 ,
input [4:0] x379 ,
input [4:0] x380 ,
input [4:0] x381 ,
input [4:0] x382 ,
input [4:0] x383 ,
input [4:0] x384 ,
input [4:0] x385 ,
input [4:0] x386 ,
input [4:0] x387 ,
input [4:0] x388 ,
input [4:0] x389 ,
input [4:0] x390 ,
input [4:0] x391 ,
input [4:0] x392 ,
input [4:0] x393 ,
input [4:0] x394 ,
input [4:0] x395 ,
input [4:0] x396 ,
input [4:0] x397 ,
input [4:0] x398 ,
input [4:0] x399 ,
input [4:0] x400 ,
input [4:0] x401 ,
input [4:0] x402 ,
input [4:0] x403 ,
input [4:0] x404 ,
input [4:0] x405 ,
input [4:0] x406 ,
input [4:0] x407 ,
input [4:0] x408 ,
input [4:0] x409 ,
input [4:0] x410 ,
input [4:0] x411 ,
input [4:0] x412 ,
input [4:0] x413 ,
input [4:0] x414 ,
input [4:0] x415 ,
input [4:0] x416 ,
input [4:0] x417 ,
input [4:0] x418 ,
input [4:0] x419 ,
input [4:0] x420 ,
input [4:0] x421 ,
input [4:0] x422 ,
input [4:0] x423 ,
input [4:0] x424 ,
input [4:0] x425 ,
input [4:0] x426 ,
input [4:0] x427 ,
input [4:0] x428 ,
input [4:0] x429 ,
input [4:0] x430 ,
input [4:0] x431 ,
input [4:0] x432 ,
input [4:0] x433 ,
input [4:0] x434 ,
input [4:0] x435 ,
input [4:0] x436 ,
input [4:0] x437 ,
input [4:0] x438 ,
input [4:0] x439 ,
input [4:0] x440 ,
input [4:0] x441 ,
input [4:0] x442 ,
input [4:0] x443 ,
input [4:0] x444 ,
input [4:0] x445 ,
input [4:0] x446 ,
input [4:0] x447 ,
input [4:0] x448 ,
input [4:0] x449 ,
input [4:0] x450 ,
input [4:0] x451 ,
input [4:0] x452 ,
input [4:0] x453 ,
input [4:0] x454 ,
input [4:0] x455 ,
input [4:0] x456 ,
input [4:0] x457 ,
input [4:0] x458 ,
input [4:0] x459 ,
input [4:0] x460 ,
input [4:0] x461 ,
input [4:0] x462 ,
input [4:0] x463 ,
input [4:0] x464 ,
input [4:0] x465 ,
input [4:0] x466 ,
input [4:0] x467 ,
input [4:0] x468 ,
input [4:0] x469 ,
input [4:0] x470 ,
input [4:0] x471 ,
input [4:0] x472 ,
input [4:0] x473 ,
input [4:0] x474 ,
input [4:0] x475 ,
input [4:0] x476 ,
input [4:0] x477 ,
input [4:0] x478 ,
input [4:0] x479 ,
input [4:0] x480 ,
input [4:0] x481 ,
input [4:0] x482 ,
input [4:0] x483 ,
input [4:0] x484 ,
input [4:0] x485 ,
input [4:0] x486 ,
input [4:0] x487 ,
input [4:0] x488 ,
input [4:0] x489 ,
input [4:0] x490 ,
input [4:0] x491 ,
input [4:0] x492 ,
input [4:0] x493 ,
input [4:0] x494 ,
input [4:0] x495 ,
output [5:0] y0 ,
output [5:0] y1 ,
output [5:0] y2 ,
output [5:0] y3 ,
output [5:0] y4 ,
output [5:0] y5 ,
output [5:0] y6 ,
output [5:0] y7 ,
output [5:0] y8 ,
output [5:0] y9 ,
output [5:0] y10 ,
output [5:0] y11 ,
output [5:0] y12 ,
output [5:0] y13 ,
output [5:0] y14 ,
output [5:0] y15 ,
output [5:0] y16 ,
output [5:0] y17 ,
output [5:0] y18 ,
output [5:0] y19 
);
wire signed[13:0] temp_y  [0:19];
assign temp_y[0] = 
+$signed( { 1'b0,x0 }  )+$signed( { 1'b0,x1 }  )+$signed( -{ 2'b0,x2 }<<<3'd1 )+$signed( { 1'b0,x3 }  )+$signed( -{ 3'b0,x6 }<<<3'd2)+$signed( { 3'b0,x7 }<<<3'd2 )+$signed( -{ 3'b0,x8 }<<<3'd2)+$signed( -{ 3'b0,x9 }<<<3'd2)+$signed( { 1'b0,x10 }  )+$signed( -{ 2'b0,x12 }<<<3'd1 )+$signed( -{ 2'b0,x13 }<<<3'd1 )+$signed( -{ 1'b0,x14 } )+$signed( -{ 1'b0,x15 } )+$signed( { 3'b0,x16 }<<<3'd2 )+$signed( { 2'b0,x17 } <<<3'd1 )+$signed( -{ 1'b0,x18 } )+$signed( { 2'b0,x19 } <<<3'd1 )+$signed( { 1'b0,x21 }  )+$signed( -{ 2'b0,x23 }<<<3'd1 )+$signed( { 2'b0,x24 } <<<3'd1 )+$signed( -{ 4'b0, x25 }<<<3'd3 )+$signed( -{ 2'b0,x26 }<<<3'd1 )+$signed( { 2'b0,x27 } <<<3'd1 )+$signed( -{ 2'b0,x28 }<<<3'd1 )+$signed( -{ 1'b0,x29 } )+$signed( -{ 3'b0,x30 }<<<3'd2)+$signed( { 1'b0,x31 }  )+$signed( { 1'b0,x32 }  )+$signed( { 1'b0,x33 }  )+$signed( { 2'b0,x34 } <<<3'd1 )+$signed( { 2'b0,x35 } <<<3'd1 )+$signed( -{ 1'b0,x36 } )+$signed( { 1'b0,x37 }  )+$signed( -{ 3'b0,x38 }<<<3'd2)+$signed( { 1'b0,x40 }  )+$signed( -{ 1'b0,x41 } )+$signed( -{ 1'b0,x42 } )+$signed( { 4'b0,x43 }<<<3'd3 )+$signed( -{ 3'b0,x44 }<<<3'd2)+$signed( { 3'b0,x45 }<<<3'd2 )+$signed( -{ 1'b0,x46 } )+$signed( -{ 2'b0,x47 }<<<3'd1 )+$signed( -{ 2'b0,x48 }<<<3'd1 )+$signed( { 2'b0,x49 } <<<3'd1 )+$signed( -{ 2'b0,x50 }<<<3'd1 )+$signed( { 2'b0,x51 } <<<3'd1 )+$signed( { 2'b0,x52 } <<<3'd1 )+$signed( { 3'b0,x53 }<<<3'd2 )+$signed( { 3'b0,x55 }<<<3'd2 )+$signed( -{ 2'b0,x56 }<<<3'd1 )+$signed( { 3'b0,x57 }<<<3'd2 )+$signed( -{ 1'b0,x59 } )+$signed( { 1'b0,x60 }  )+$signed( -{ 1'b0,x61 } )+$signed( -{ 3'b0,x62 }<<<3'd2)+$signed( { 3'b0,x63 }<<<3'd2 )+$signed( { 2'b0,x64 } <<<3'd1 )+$signed( { 1'b0,x65 }  )+$signed( { 1'b0,x66 }  )+$signed( { 1'b0,x67 }  )+$signed( -{ 2'b0,x68 }<<<3'd1 )+$signed( { 2'b0,x69 } <<<3'd1 )+$signed( -{ 1'b0,x70 } )+$signed( { 3'b0,x71 }<<<3'd2 )+$signed( -{ 3'b0,x72 }<<<3'd2)+$signed( { 3'b0,x73 }<<<3'd2 )+$signed( { 2'b0,x74 } <<<3'd1 )+$signed( { 2'b0,x75 } <<<3'd1 )+$signed( { 1'b0,x76 }  )+$signed( { 2'b0,x78 } <<<3'd1 )+$signed( -{ 2'b0,x79 }<<<3'd1 )+$signed( -{ 4'b0, x80 }<<<3'd3 )+$signed( { 1'b0,x81 }  )+$signed( -{ 1'b0,x82 } )+$signed( { 3'b0,x84 }<<<3'd2 )+$signed( -{ 1'b0,x85 } )+$signed( -{ 3'b0,x86 }<<<3'd2)+$signed( { 3'b0,x88 }<<<3'd2 )+$signed( { 2'b0,x89 } <<<3'd1 )+$signed( -{ 1'b0,x91 } )+$signed( -{ 3'b0,x92 }<<<3'd2)+$signed( -{ 2'b0,x93 }<<<3'd1 )+$signed( -{ 2'b0,x94 }<<<3'd1 )+$signed( -{ 2'b0,x95 }<<<3'd1 )+$signed( { 3'b0,x96 }<<<3'd2 )+$signed( { 2'b0,x97 } <<<3'd1 )+$signed( { 5'b0,x98  }<<<3'd4 )+$signed( -{ 3'b0,x100 }<<<3'd2)+$signed( -{ 4'b0, x101 }<<<3'd3 )+$signed( -{ 2'b0,x102 }<<<3'd1 )+$signed( { 3'b0,x104 }<<<3'd2 )+$signed( -{ 2'b0,x105 }<<<3'd1 )+$signed( -{ 3'b0,x107 }<<<3'd2)+$signed( -{ 1'b0,x108 } )+$signed( -{ 3'b0,x109 }<<<3'd2)+$signed( -{ 1'b0,x111 } )+$signed( { 1'b0,x112 }  )+$signed( -{ 3'b0,x113 }<<<3'd2)+$signed( -{ 1'b0,x114 } )+$signed( { 5'b0,x116  }<<<3'd4 )+$signed( { 3'b0,x117 }<<<3'd2 )+$signed( { 2'b0,x118 } <<<3'd1 )+$signed( -{ 4'b0, x119 }<<<3'd3 )+$signed( -{ 3'b0,x120 }<<<3'd2)+$signed( -{ 2'b0,x121 }<<<3'd1 )+$signed( { 1'b0,x122 }  )+$signed( { 1'b0,x124 }  )+$signed( -{ 4'b0, x125 }<<<3'd3 )+$signed( -{ 1'b0,x126 } )+$signed( { 2'b0,x127 } <<<3'd1 )+$signed( -{ 2'b0,x128 }<<<3'd1 )+$signed( -{ 3'b0,x129 }<<<3'd2)+$signed( { 2'b0,x130 } <<<3'd1 )+$signed( { 3'b0,x131 }<<<3'd2 )+$signed( { 3'b0,x132 }<<<3'd2 )+$signed( { 3'b0,x133 }<<<3'd2 )+$signed( -{ 4'b0, x134 }<<<3'd3 )+$signed( { 1'b0,x135 }  )+$signed( { 2'b0,x136 } <<<3'd1 )+$signed( { 3'b0,x137 }<<<3'd2 )+$signed( { 3'b0,x139 }<<<3'd2 )+$signed( -{ 3'b0,x140 }<<<3'd2)+$signed( { 3'b0,x142 }<<<3'd2 )+$signed( { 1'b0,x143 }  )+$signed( -{ 2'b0,x144 }<<<3'd1 )+$signed( { 3'b0,x145 }<<<3'd2 )+$signed( { 1'b0,x147 }  )+$signed( -{ 1'b0,x148 } )+$signed( -{ 2'b0,x149 }<<<3'd1 )+$signed( { 2'b0,x150 } <<<3'd1 )+$signed( { 1'b0,x151 }  )+$signed( -{ 3'b0,x152 }<<<3'd2)+$signed( -{ 1'b0,x154 } )+$signed( { 1'b0,x155 }  )+$signed( -{ 1'b0,x156 } )+$signed( -{ 3'b0,x157 }<<<3'd2)+$signed( -{ 2'b0,x158 }<<<3'd1 )+$signed( -{ 2'b0,x159 }<<<3'd1 )+$signed( { 3'b0,x160 }<<<3'd2 )+$signed( { 2'b0,x161 } <<<3'd1 )+$signed( -{ 2'b0,x162 }<<<3'd1 )+$signed( -{ 2'b0,x163 }<<<3'd1 )+$signed( -{ 1'b0,x164 } )+$signed( -{ 3'b0,x165 }<<<3'd2)+$signed( -{ 2'b0,x166 }<<<3'd1 )+$signed( -{ 3'b0,x167 }<<<3'd2)+$signed( { 1'b0,x168 }  )+$signed( -{ 2'b0,x169 }<<<3'd1 )+$signed( { 4'b0,x170 }<<<3'd3 )+$signed( -{ 3'b0,x171 }<<<3'd2)+$signed( { 2'b0,x172 } <<<3'd1 )+$signed( { 2'b0,x174 } <<<3'd1 )+$signed( -{ 1'b0,x175 } )+$signed( -{ 2'b0,x176 }<<<3'd1 )+$signed( { 1'b0,x177 }  )+$signed( { 2'b0,x178 } <<<3'd1 )+$signed( -{ 1'b0,x179 } )+$signed( -{ 3'b0,x180 }<<<3'd2)+$signed( -{ 1'b0,x181 } )+$signed( { 2'b0,x182 } <<<3'd1 )+$signed( -{ 3'b0,x183 }<<<3'd2)+$signed( -{ 2'b0,x184 }<<<3'd1 )+$signed( -{ 1'b0,x185 } )+$signed( { 3'b0,x186 }<<<3'd2 )+$signed( { 3'b0,x187 }<<<3'd2 )+$signed( { 4'b0,x188 }<<<3'd3 )+$signed( -{ 2'b0,x189 }<<<3'd1 )+$signed( { 2'b0,x190 } <<<3'd1 )+$signed( -{ 2'b0,x191 }<<<3'd1 )+$signed( -{ 2'b0,x193 }<<<3'd1 )+$signed( -{ 1'b0,x194 } )+$signed( -{ 1'b0,x197 } )+$signed( { 2'b0,x198 } <<<3'd1 )+$signed( { 1'b0,x199 }  )+$signed( -{ 1'b0,x200 } )+$signed( -{ 2'b0,x201 }<<<3'd1 )+$signed( -{ 1'b0,x202 } )+$signed( -{ 2'b0,x203 }<<<3'd1 )+$signed( { 2'b0,x204 } <<<3'd1 )+$signed( -{ 3'b0,x206 }<<<3'd2)+$signed( -{ 2'b0,x207 }<<<3'd1 )+$signed( { 3'b0,x208 }<<<3'd2 )+$signed( { 1'b0,x209 }  )+$signed( -{ 3'b0,x210 }<<<3'd2)+$signed( -{ 2'b0,x211 }<<<3'd1 )+$signed( { 3'b0,x212 }<<<3'd2 )+$signed( { 2'b0,x213 } <<<3'd1 )+$signed( { 2'b0,x216 } <<<3'd1 )+$signed( { 4'b0,x217 }<<<3'd3 )+$signed( { 2'b0,x219 } <<<3'd1 )+$signed( { 3'b0,x221 }<<<3'd2 )+$signed( { 2'b0,x222 } <<<3'd1 )+$signed( { 2'b0,x223 } <<<3'd1 )+$signed( -{ 3'b0,x224 }<<<3'd2)+$signed( -{ 3'b0,x225 }<<<3'd2)+$signed( { 3'b0,x226 }<<<3'd2 )+$signed( { 1'b0,x227 }  )+$signed( -{ 1'b0,x228 } )+$signed( -{ 2'b0,x229 }<<<3'd1 )+$signed( -{ 3'b0,x230 }<<<3'd2)+$signed( -{ 1'b0,x232 } )+$signed( { 2'b0,x233 } <<<3'd1 )+$signed( { 3'b0,x235 }<<<3'd2 )+$signed( { 1'b0,x236 }  )+$signed( { 3'b0,x237 }<<<3'd2 )+$signed( { 2'b0,x238 } <<<3'd1 )+$signed( -{ 1'b0,x239 } )+$signed( -{ 1'b0,x240 } )+$signed( -{ 1'b0,x241 } )+$signed( -{ 3'b0,x242 }<<<3'd2)+$signed( -{ 3'b0,x243 }<<<3'd2)+$signed( { 2'b0,x244 } <<<3'd1 )+$signed( { 2'b0,x245 } <<<3'd1 )+$signed( -{ 3'b0,x246 }<<<3'd2)+$signed( -{ 3'b0,x247 }<<<3'd2)+$signed( -{ 2'b0,x248 }<<<3'd1 )+$signed( -{ 3'b0,x249 }<<<3'd2)+$signed( -{ 2'b0,x250 }<<<3'd1 )+$signed( { 3'b0,x251 }<<<3'd2 )+$signed( { 2'b0,x253 } <<<3'd1 )+$signed( { 2'b0,x254 } <<<3'd1 )+$signed( { 3'b0,x255 }<<<3'd2 )+$signed( { 1'b0,x256 }  )+$signed( { 2'b0,x257 } <<<3'd1 )+$signed( { 3'b0,x258 }<<<3'd2 )+$signed( -{ 2'b0,x259 }<<<3'd1 )+$signed( -{ 1'b0,x260 } )+$signed( -{ 4'b0, x261 }<<<3'd3 )+$signed( { 3'b0,x262 }<<<3'd2 )+$signed( { 3'b0,x263 }<<<3'd2 )+$signed( { 1'b0,x264 }  )+$signed( -{ 4'b0, x265 }<<<3'd3 )+$signed( { 2'b0,x266 } <<<3'd1 )+$signed( -{ 2'b0,x267 }<<<3'd1 )+$signed( -{ 2'b0,x268 }<<<3'd1 )+$signed( { 1'b0,x269 }  )+$signed( { 2'b0,x270 } <<<3'd1 )+$signed( { 1'b0,x271 }  )+$signed( -{ 2'b0,x272 }<<<3'd1 )+$signed( { 4'b0,x273 }<<<3'd3 )+$signed( -{ 2'b0,x274 }<<<3'd1 )+$signed( { 1'b0,x275 }  )+$signed( { 3'b0,x276 }<<<3'd2 )+$signed( -{ 3'b0,x277 }<<<3'd2)+$signed( -{ 3'b0,x278 }<<<3'd2)+$signed( -{ 3'b0,x279 }<<<3'd2)+$signed( { 3'b0,x280 }<<<3'd2 )+$signed( -{ 2'b0,x281 }<<<3'd1 )+$signed( -{ 1'b0,x282 } )+$signed( -{ 2'b0,x283 }<<<3'd1 )+$signed( -{ 2'b0,x284 }<<<3'd1 )+$signed( -{ 3'b0,x286 }<<<3'd2)+$signed( { 2'b0,x287 } <<<3'd1 )+$signed( { 3'b0,x288 }<<<3'd2 )+$signed( { 1'b0,x289 }  )+$signed( -{ 3'b0,x290 }<<<3'd2)+$signed( { 2'b0,x291 } <<<3'd1 )+$signed( -{ 1'b0,x292 } )+$signed( -{ 2'b0,x294 }<<<3'd1 )+$signed( -{ 1'b0,x295 } )+$signed( -{ 2'b0,x297 }<<<3'd1 )+$signed( -{ 2'b0,x298 }<<<3'd1 )+$signed( { 2'b0,x299 } <<<3'd1 )+$signed( { 2'b0,x300 } <<<3'd1 )+$signed( -{ 2'b0,x301 }<<<3'd1 )+$signed( { 1'b0,x303 }  )+$signed( { 1'b0,x304 }  )+$signed( -{ 1'b0,x305 } )+$signed( -{ 3'b0,x306 }<<<3'd2)+$signed( -{ 2'b0,x307 }<<<3'd1 )+$signed( { 3'b0,x308 }<<<3'd2 )+$signed( -{ 3'b0,x309 }<<<3'd2)+$signed( { 3'b0,x311 }<<<3'd2 )+$signed( { 3'b0,x312 }<<<3'd2 )+$signed( { 2'b0,x313 } <<<3'd1 )+$signed( -{ 3'b0,x315 }<<<3'd2)+$signed( -{ 1'b0,x316 } )+$signed( -{ 3'b0,x317 }<<<3'd2)+$signed( -{ 2'b0,x318 }<<<3'd1 )+$signed( -{ 3'b0,x319 }<<<3'd2)+$signed( -{ 1'b0,x320 } )+$signed( { 1'b0,x321 }  )+$signed( -{ 1'b0,x322 } )+$signed( { 2'b0,x323 } <<<3'd1 )+$signed( -{ 2'b0,x324 }<<<3'd1 )+$signed( { 2'b0,x325 } <<<3'd1 )+$signed( { 1'b0,x326 }  )+$signed( { 2'b0,x327 } <<<3'd1 )+$signed( { 1'b0,x328 }  )+$signed( { 1'b0,x329 }  )+$signed( { 2'b0,x330 } <<<3'd1 )+$signed( { 3'b0,x331 }<<<3'd2 )+$signed( { 1'b0,x332 }  )+$signed( { 2'b0,x334 } <<<3'd1 )+$signed( { 1'b0,x335 }  )+$signed( -{ 3'b0,x336 }<<<3'd2)+$signed( { 2'b0,x338 } <<<3'd1 )+$signed( -{ 2'b0,x339 }<<<3'd1 )+$signed( -{ 3'b0,x340 }<<<3'd2)+$signed( { 3'b0,x341 }<<<3'd2 )+$signed( -{ 1'b0,x342 } )+$signed( { 3'b0,x343 }<<<3'd2 )+$signed( -{ 2'b0,x344 }<<<3'd1 )+$signed( -{ 2'b0,x345 }<<<3'd1 )+$signed( { 2'b0,x346 } <<<3'd1 )+$signed( { 1'b0,x347 }  )+$signed( { 1'b0,x348 }  )+$signed( { 2'b0,x349 } <<<3'd1 )+$signed( { 1'b0,x351 }  )+$signed( -{ 3'b0,x353 }<<<3'd2)+$signed( -{ 3'b0,x355 }<<<3'd2)+$signed( -{ 1'b0,x357 } )+$signed( -{ 2'b0,x359 }<<<3'd1 )+$signed( { 2'b0,x360 } <<<3'd1 )+$signed( { 2'b0,x361 } <<<3'd1 )+$signed( { 5'b0,x362  }<<<3'd4 )+$signed( -{ 1'b0,x363 } )+$signed( { 2'b0,x364 } <<<3'd1 )+$signed( { 3'b0,x365 }<<<3'd2 )+$signed( { 2'b0,x366 } <<<3'd1 )+$signed( { 3'b0,x367 }<<<3'd2 )+$signed( -{ 1'b0,x368 } )+$signed( { 3'b0,x370 }<<<3'd2 )+$signed( -{ 3'b0,x372 }<<<3'd2)+$signed( -{ 3'b0,x374 }<<<3'd2)+$signed( { 4'b0,x375 }<<<3'd3 )+$signed( -{ 2'b0,x376 }<<<3'd1 )+$signed( -{ 3'b0,x377 }<<<3'd2)+$signed( { 3'b0,x379 }<<<3'd2 )+$signed( { 3'b0,x380 }<<<3'd2 )+$signed( -{ 2'b0,x381 }<<<3'd1 )+$signed( -{ 3'b0,x382 }<<<3'd2)+$signed( -{ 4'b0, x383 }<<<3'd3 )+$signed( -{ 1'b0,x385 } )+$signed( { 2'b0,x386 } <<<3'd1 )+$signed( -{ 2'b0,x387 }<<<3'd1 )+$signed( -{ 4'b0, x388 }<<<3'd3 )+$signed( -{ 3'b0,x390 }<<<3'd2)+$signed( -{ 2'b0,x391 }<<<3'd1 )+$signed( -{ 3'b0,x392 }<<<3'd2)+$signed( { 1'b0,x393 }  )+$signed( { 2'b0,x394 } <<<3'd1 )+$signed( { 3'b0,x395 }<<<3'd2 )+$signed( { 3'b0,x396 }<<<3'd2 )+$signed( -{ 3'b0,x397 }<<<3'd2)+$signed( { 1'b0,x398 }  )+$signed( { 1'b0,x399 }  )+$signed( { 3'b0,x400 }<<<3'd2 )+$signed( -{ 2'b0,x401 }<<<3'd1 )+$signed( { 1'b0,x402 }  )+$signed( { 3'b0,x403 }<<<3'd2 )+$signed( { 3'b0,x406 }<<<3'd2 )+$signed( -{ 2'b0,x407 }<<<3'd1 )+$signed( -{ 1'b0,x408 } )+$signed( -{ 2'b0,x409 }<<<3'd1 )+$signed( -{ 2'b0,x411 }<<<3'd1 )+$signed( { 2'b0,x412 } <<<3'd1 )+$signed( { 2'b0,x413 } <<<3'd1 )+$signed( { 1'b0,x414 }  )+$signed( -{ 1'b0,x417 } )+$signed( -{ 3'b0,x418 }<<<3'd2)+$signed( { 2'b0,x419 } <<<3'd1 )+$signed( { 1'b0,x420 }  )+$signed( -{ 3'b0,x422 }<<<3'd2)+$signed( -{ 2'b0,x423 }<<<3'd1 )+$signed( { 3'b0,x426 }<<<3'd2 )+$signed( -{ 1'b0,x427 } )+$signed( { 1'b0,x429 }  )+$signed( -{ 2'b0,x430 }<<<3'd1 )+$signed( -{ 3'b0,x431 }<<<3'd2)+$signed( { 3'b0,x432 }<<<3'd2 )+$signed( -{ 1'b0,x433 } )+$signed( -{ 3'b0,x434 }<<<3'd2)+$signed( -{ 3'b0,x435 }<<<3'd2)+$signed( { 2'b0,x436 } <<<3'd1 )+$signed( -{ 1'b0,x437 } )+$signed( { 3'b0,x438 }<<<3'd2 )+$signed( -{ 3'b0,x439 }<<<3'd2)+$signed( -{ 3'b0,x440 }<<<3'd2)+$signed( -{ 1'b0,x441 } )+$signed( -{ 2'b0,x442 }<<<3'd1 )+$signed( -{ 1'b0,x443 } )+$signed( -{ 1'b0,x444 } )+$signed( { 3'b0,x445 }<<<3'd2 )+$signed( { 2'b0,x446 } <<<3'd1 )+$signed( -{ 1'b0,x447 } )+$signed( { 1'b0,x448 }  )+$signed( -{ 2'b0,x449 }<<<3'd1 )+$signed( -{ 3'b0,x452 }<<<3'd2)+$signed( -{ 4'b0, x453 }<<<3'd3 )+$signed( -{ 2'b0,x454 }<<<3'd1 )+$signed( { 4'b0,x455 }<<<3'd3 )+$signed( { 2'b0,x456 } <<<3'd1 )+$signed( -{ 1'b0,x457 } )+$signed( { 3'b0,x458 }<<<3'd2 )+$signed( { 1'b0,x459 }  )+$signed( { 2'b0,x460 } <<<3'd1 )+$signed( { 2'b0,x461 } <<<3'd1 )+$signed( -{ 2'b0,x462 }<<<3'd1 )+$signed( -{ 1'b0,x463 } )+$signed( { 3'b0,x464 }<<<3'd2 )+$signed( -{ 1'b0,x465 } )+$signed( -{ 3'b0,x466 }<<<3'd2)+$signed( -{ 3'b0,x467 }<<<3'd2)+$signed( { 4'b0,x468 }<<<3'd3 )+$signed( -{ 3'b0,x469 }<<<3'd2)+$signed( { 1'b0,x470 }  )+$signed( -{ 1'b0,x471 } )+$signed( -{ 2'b0,x473 }<<<3'd1 )+$signed( -{ 3'b0,x474 }<<<3'd2)+$signed( { 2'b0,x475 } <<<3'd1 )+$signed( -{ 2'b0,x476 }<<<3'd1 )+$signed( { 3'b0,x477 }<<<3'd2 )+$signed( -{ 3'b0,x479 }<<<3'd2)+$signed( -{ 2'b0,x480 }<<<3'd1 )+$signed( { 2'b0,x481 } <<<3'd1 )+$signed( -{ 3'b0,x482 }<<<3'd2)+$signed( { 2'b0,x483 } <<<3'd1 )+$signed( -{ 2'b0,x484 }<<<3'd1 )+$signed( { 2'b0,x485 } <<<3'd1 )+$signed( -{ 3'b0,x486 }<<<3'd2)+$signed( -{ 4'b0, x487 }<<<3'd3 )+$signed( -{ 3'b0,x488 }<<<3'd2)+$signed( -{ 2'b0,x489 }<<<3'd1 )+$signed( { 1'b0,x490 }  )+$signed( -{ 1'b0,x491 } )+$signed( -{ 1'b0,x492 } )+$signed( -{ 3'b0,x493 }<<<3'd2)+$signed( { 2'b0,x495 } <<<3'd1 )-$signed(13'd16);
assign y0=temp_y[0][13] ==1'b1 ? 6'd0 :  
    temp_y[0][10] ==1'b1 ? 6'd63 : 
    temp_y[0][3]==1'b1 ? temp_y[0][9:4]+1'b1 : temp_y[0][9:4];
assign temp_y[1] = 
+$signed( -{ 3'b0,x1 }<<<3'd2)+$signed( -{ 2'b0,x2 }<<<3'd1 )+$signed( -{ 4'b0, x3 }<<<3'd3 )+$signed( -{ 2'b0,x4 }<<<3'd1 )+$signed( -{ 2'b0,x5 }<<<3'd1 )+$signed( { 5'b0,x7  }<<<3'd4 )+$signed( -{ 2'b0,x8 }<<<3'd1 )+$signed( -{ 2'b0,x9 }<<<3'd1 )+$signed( { 3'b0,x10 }<<<3'd2 )+$signed( -{ 4'b0, x11 }<<<3'd3 )+$signed( -{ 3'b0,x12 }<<<3'd2)+$signed( -{ 2'b0,x13 }<<<3'd1 )+$signed( -{ 2'b0,x14 }<<<3'd1 )+$signed( { 4'b0,x15 }<<<3'd3 )+$signed( -{ 1'b0,x16 } )+$signed( -{ 4'b0, x17 }<<<3'd3 )+$signed( -{ 3'b0,x18 }<<<3'd2)+$signed( -{ 1'b0,x19 } )+$signed( -{ 2'b0,x20 }<<<3'd1 )+$signed( -{ 3'b0,x21 }<<<3'd2)+$signed( { 3'b0,x22 }<<<3'd2 )+$signed( -{ 3'b0,x23 }<<<3'd2)+$signed( { 4'b0,x25 }<<<3'd3 )+$signed( { 1'b0,x26 }  )+$signed( -{ 1'b0,x27 } )+$signed( { 3'b0,x28 }<<<3'd2 )+$signed( -{ 3'b0,x29 }<<<3'd2)+$signed( -{ 3'b0,x30 }<<<3'd2)+$signed( -{ 2'b0,x31 }<<<3'd1 )+$signed( -{ 2'b0,x33 }<<<3'd1 )+$signed( -{ 2'b0,x34 }<<<3'd1 )+$signed( -{ 3'b0,x35 }<<<3'd2)+$signed( { 1'b0,x37 }  )+$signed( -{ 1'b0,x38 } )+$signed( -{ 3'b0,x39 }<<<3'd2)+$signed( { 1'b0,x40 }  )+$signed( -{ 3'b0,x41 }<<<3'd2)+$signed( { 1'b0,x42 }  )+$signed( { 4'b0,x43 }<<<3'd3 )+$signed( -{ 1'b0,x44 } )+$signed( -{ 1'b0,x45 } )+$signed( { 2'b0,x46 } <<<3'd1 )+$signed( -{ 3'b0,x47 }<<<3'd2)+$signed( -{ 3'b0,x48 }<<<3'd2)+$signed( -{ 3'b0,x49 }<<<3'd2)+$signed( { 3'b0,x50 }<<<3'd2 )+$signed( { 1'b0,x51 }  )+$signed( -{ 1'b0,x52 } )+$signed( -{ 4'b0, x53 }<<<3'd3 )+$signed( -{ 2'b0,x54 }<<<3'd1 )+$signed( { 2'b0,x55 } <<<3'd1 )+$signed( -{ 3'b0,x56 }<<<3'd2)+$signed( -{ 2'b0,x57 }<<<3'd1 )+$signed( -{ 3'b0,x58 }<<<3'd2)+$signed( -{ 3'b0,x59 }<<<3'd2)+$signed( -{ 1'b0,x61 } )+$signed( { 2'b0,x63 } <<<3'd1 )+$signed( { 3'b0,x64 }<<<3'd2 )+$signed( -{ 1'b0,x65 } )+$signed( { 1'b0,x68 }  )+$signed( -{ 3'b0,x69 }<<<3'd2)+$signed( -{ 1'b0,x70 } )+$signed( -{ 4'b0, x71 }<<<3'd3 )+$signed( { 1'b0,x72 }  )+$signed( -{ 3'b0,x73 }<<<3'd2)+$signed( { 2'b0,x74 } <<<3'd1 )+$signed( -{ 3'b0,x75 }<<<3'd2)+$signed( -{ 3'b0,x77 }<<<3'd2)+$signed( -{ 1'b0,x79 } )+$signed( -{ 2'b0,x80 }<<<3'd1 )+$signed( -{ 1'b0,x81 } )+$signed( { 2'b0,x82 } <<<3'd1 )+$signed( { 2'b0,x83 } <<<3'd1 )+$signed( -{ 2'b0,x84 }<<<3'd1 )+$signed( -{ 2'b0,x85 }<<<3'd1 )+$signed( -{ 1'b0,x86 } )+$signed( -{ 2'b0,x88 }<<<3'd1 )+$signed( -{ 3'b0,x89 }<<<3'd2)+$signed( -{ 3'b0,x91 }<<<3'd2)+$signed( -{ 2'b0,x92 }<<<3'd1 )+$signed( -{ 4'b0, x93 }<<<3'd3 )+$signed( -{ 2'b0,x94 }<<<3'd1 )+$signed( -{ 3'b0,x95 }<<<3'd2)+$signed( -{ 2'b0,x96 }<<<3'd1 )+$signed( { 2'b0,x97 } <<<3'd1 )+$signed( -{ 1'b0,x100 } )+$signed( { 3'b0,x101 }<<<3'd2 )+$signed( -{ 2'b0,x102 }<<<3'd1 )+$signed( -{ 4'b0, x104 }<<<3'd3 )+$signed( { 2'b0,x105 } <<<3'd1 )+$signed( { 2'b0,x106 } <<<3'd1 )+$signed( -{ 3'b0,x107 }<<<3'd2)+$signed( { 3'b0,x108 }<<<3'd2 )+$signed( -{ 3'b0,x110 }<<<3'd2)+$signed( -{ 3'b0,x111 }<<<3'd2)+$signed( -{ 2'b0,x112 }<<<3'd1 )+$signed( -{ 1'b0,x113 } )+$signed( -{ 2'b0,x114 }<<<3'd1 )+$signed( { 3'b0,x115 }<<<3'd2 )+$signed( -{ 1'b0,x116 } )+$signed( -{ 2'b0,x117 }<<<3'd1 )+$signed( -{ 3'b0,x118 }<<<3'd2)+$signed( { 2'b0,x119 } <<<3'd1 )+$signed( { 1'b0,x120 }  )+$signed( { 1'b0,x121 }  )+$signed( -{ 4'b0, x122 }<<<3'd3 )+$signed( { 3'b0,x123 }<<<3'd2 )+$signed( { 1'b0,x124 }  )+$signed( -{ 1'b0,x125 } )+$signed( { 2'b0,x126 } <<<3'd1 )+$signed( -{ 2'b0,x127 }<<<3'd1 )+$signed( -{ 2'b0,x128 }<<<3'd1 )+$signed( -{ 4'b0, x129 }<<<3'd3 )+$signed( { 1'b0,x130 }  )+$signed( { 3'b0,x132 }<<<3'd2 )+$signed( { 3'b0,x133 }<<<3'd2 )+$signed( -{ 3'b0,x134 }<<<3'd2)+$signed( { 3'b0,x136 }<<<3'd2 )+$signed( -{ 3'b0,x137 }<<<3'd2)+$signed( -{ 1'b0,x138 } )+$signed( { 2'b0,x139 } <<<3'd1 )+$signed( -{ 3'b0,x140 }<<<3'd2)+$signed( -{ 3'b0,x141 }<<<3'd2)+$signed( { 3'b0,x142 }<<<3'd2 )+$signed( -{ 1'b0,x143 } )+$signed( { 1'b0,x144 }  )+$signed( { 2'b0,x145 } <<<3'd1 )+$signed( -{ 3'b0,x146 }<<<3'd2)+$signed( { 3'b0,x147 }<<<3'd2 )+$signed( { 2'b0,x148 } <<<3'd1 )+$signed( -{ 1'b0,x149 } )+$signed( { 2'b0,x152 } <<<3'd1 )+$signed( -{ 2'b0,x153 }<<<3'd1 )+$signed( -{ 1'b0,x154 } )+$signed( { 3'b0,x155 }<<<3'd2 )+$signed( { 2'b0,x156 } <<<3'd1 )+$signed( { 2'b0,x157 } <<<3'd1 )+$signed( { 2'b0,x158 } <<<3'd1 )+$signed( -{ 2'b0,x160 }<<<3'd1 )+$signed( { 1'b0,x161 }  )+$signed( -{ 2'b0,x162 }<<<3'd1 )+$signed( { 2'b0,x163 } <<<3'd1 )+$signed( { 2'b0,x164 } <<<3'd1 )+$signed( -{ 3'b0,x165 }<<<3'd2)+$signed( -{ 2'b0,x166 }<<<3'd1 )+$signed( { 3'b0,x167 }<<<3'd2 )+$signed( -{ 2'b0,x169 }<<<3'd1 )+$signed( { 2'b0,x170 } <<<3'd1 )+$signed( { 2'b0,x171 } <<<3'd1 )+$signed( { 1'b0,x172 }  )+$signed( { 3'b0,x173 }<<<3'd2 )+$signed( -{ 2'b0,x176 }<<<3'd1 )+$signed( { 3'b0,x178 }<<<3'd2 )+$signed( -{ 2'b0,x179 }<<<3'd1 )+$signed( { 2'b0,x180 } <<<3'd1 )+$signed( { 3'b0,x181 }<<<3'd2 )+$signed( -{ 1'b0,x182 } )+$signed( -{ 3'b0,x183 }<<<3'd2)+$signed( -{ 3'b0,x184 }<<<3'd2)+$signed( { 1'b0,x185 }  )+$signed( -{ 1'b0,x187 } )+$signed( { 3'b0,x188 }<<<3'd2 )+$signed( -{ 2'b0,x189 }<<<3'd1 )+$signed( -{ 2'b0,x190 }<<<3'd1 )+$signed( { 4'b0,x191 }<<<3'd3 )+$signed( { 2'b0,x192 } <<<3'd1 )+$signed( { 2'b0,x193 } <<<3'd1 )+$signed( -{ 2'b0,x194 }<<<3'd1 )+$signed( { 3'b0,x196 }<<<3'd2 )+$signed( -{ 3'b0,x197 }<<<3'd2)+$signed( { 1'b0,x198 }  )+$signed( { 2'b0,x199 } <<<3'd1 )+$signed( -{ 2'b0,x200 }<<<3'd1 )+$signed( -{ 2'b0,x201 }<<<3'd1 )+$signed( -{ 1'b0,x202 } )+$signed( { 1'b0,x204 }  )+$signed( { 3'b0,x205 }<<<3'd2 )+$signed( -{ 2'b0,x206 }<<<3'd1 )+$signed( { 2'b0,x207 } <<<3'd1 )+$signed( -{ 1'b0,x208 } )+$signed( { 3'b0,x209 }<<<3'd2 )+$signed( -{ 2'b0,x210 }<<<3'd1 )+$signed( -{ 3'b0,x211 }<<<3'd2)+$signed( { 1'b0,x213 }  )+$signed( -{ 2'b0,x216 }<<<3'd1 )+$signed( { 3'b0,x217 }<<<3'd2 )+$signed( { 1'b0,x218 }  )+$signed( -{ 1'b0,x220 } )+$signed( { 3'b0,x221 }<<<3'd2 )+$signed( -{ 1'b0,x223 } )+$signed( { 2'b0,x224 } <<<3'd1 )+$signed( -{ 1'b0,x225 } )+$signed( -{ 3'b0,x226 }<<<3'd2)+$signed( { 3'b0,x227 }<<<3'd2 )+$signed( { 2'b0,x228 } <<<3'd1 )+$signed( { 3'b0,x229 }<<<3'd2 )+$signed( { 2'b0,x230 } <<<3'd1 )+$signed( -{ 2'b0,x231 }<<<3'd1 )+$signed( { 1'b0,x232 }  )+$signed( { 3'b0,x233 }<<<3'd2 )+$signed( -{ 1'b0,x234 } )+$signed( { 3'b0,x235 }<<<3'd2 )+$signed( { 3'b0,x236 }<<<3'd2 )+$signed( -{ 3'b0,x237 }<<<3'd2)+$signed( -{ 4'b0, x238 }<<<3'd3 )+$signed( { 2'b0,x239 } <<<3'd1 )+$signed( { 2'b0,x240 } <<<3'd1 )+$signed( { 2'b0,x241 } <<<3'd1 )+$signed( { 2'b0,x242 } <<<3'd1 )+$signed( -{ 2'b0,x243 }<<<3'd1 )+$signed( -{ 3'b0,x244 }<<<3'd2)+$signed( { 2'b0,x245 } <<<3'd1 )+$signed( { 1'b0,x246 }  )+$signed( { 1'b0,x247 }  )+$signed( { 3'b0,x248 }<<<3'd2 )+$signed( -{ 2'b0,x249 }<<<3'd1 )+$signed( { 2'b0,x250 } <<<3'd1 )+$signed( -{ 1'b0,x251 } )+$signed( { 1'b0,x252 }  )+$signed( { 4'b0,x253 }<<<3'd3 )+$signed( -{ 2'b0,x254 }<<<3'd1 )+$signed( -{ 2'b0,x255 }<<<3'd1 )+$signed( -{ 3'b0,x256 }<<<3'd2)+$signed( { 2'b0,x257 } <<<3'd1 )+$signed( { 3'b0,x258 }<<<3'd2 )+$signed( { 1'b0,x259 }  )+$signed( { 2'b0,x260 } <<<3'd1 )+$signed( { 2'b0,x261 } <<<3'd1 )+$signed( -{ 3'b0,x262 }<<<3'd2)+$signed( { 3'b0,x263 }<<<3'd2 )+$signed( -{ 2'b0,x264 }<<<3'd1 )+$signed( -{ 2'b0,x265 }<<<3'd1 )+$signed( { 3'b0,x266 }<<<3'd2 )+$signed( -{ 3'b0,x267 }<<<3'd2)+$signed( -{ 1'b0,x268 } )+$signed( { 2'b0,x269 } <<<3'd1 )+$signed( { 3'b0,x270 }<<<3'd2 )+$signed( { 2'b0,x272 } <<<3'd1 )+$signed( -{ 2'b0,x273 }<<<3'd1 )+$signed( -{ 1'b0,x276 } )+$signed( { 2'b0,x278 } <<<3'd1 )+$signed( -{ 3'b0,x279 }<<<3'd2)+$signed( { 3'b0,x281 }<<<3'd2 )+$signed( -{ 2'b0,x282 }<<<3'd1 )+$signed( { 1'b0,x283 }  )+$signed( { 3'b0,x284 }<<<3'd2 )+$signed( { 2'b0,x285 } <<<3'd1 )+$signed( -{ 3'b0,x286 }<<<3'd2)+$signed( { 3'b0,x287 }<<<3'd2 )+$signed( -{ 2'b0,x288 }<<<3'd1 )+$signed( { 2'b0,x289 } <<<3'd1 )+$signed( { 2'b0,x290 } <<<3'd1 )+$signed( -{ 2'b0,x291 }<<<3'd1 )+$signed( -{ 2'b0,x292 }<<<3'd1 )+$signed( -{ 4'b0, x293 }<<<3'd3 )+$signed( -{ 1'b0,x294 } )+$signed( { 3'b0,x295 }<<<3'd2 )+$signed( { 3'b0,x296 }<<<3'd2 )+$signed( { 1'b0,x298 }  )+$signed( -{ 5'b0,x299 }<<<3'd4 )+$signed( { 3'b0,x300 }<<<3'd2 )+$signed( -{ 2'b0,x301 }<<<3'd1 )+$signed( -{ 2'b0,x302 }<<<3'd1 )+$signed( { 2'b0,x303 } <<<3'd1 )+$signed( -{ 4'b0, x304 }<<<3'd3 )+$signed( { 3'b0,x305 }<<<3'd2 )+$signed( -{ 3'b0,x306 }<<<3'd2)+$signed( -{ 3'b0,x307 }<<<3'd2)+$signed( { 3'b0,x309 }<<<3'd2 )+$signed( -{ 2'b0,x310 }<<<3'd1 )+$signed( -{ 3'b0,x311 }<<<3'd2)+$signed( { 2'b0,x312 } <<<3'd1 )+$signed( { 3'b0,x313 }<<<3'd2 )+$signed( -{ 2'b0,x314 }<<<3'd1 )+$signed( -{ 2'b0,x315 }<<<3'd1 )+$signed( -{ 3'b0,x316 }<<<3'd2)+$signed( -{ 2'b0,x317 }<<<3'd1 )+$signed( { 3'b0,x318 }<<<3'd2 )+$signed( { 1'b0,x321 }  )+$signed( { 2'b0,x322 } <<<3'd1 )+$signed( { 2'b0,x323 } <<<3'd1 )+$signed( -{ 3'b0,x324 }<<<3'd2)+$signed( -{ 2'b0,x325 }<<<3'd1 )+$signed( { 3'b0,x326 }<<<3'd2 )+$signed( { 1'b0,x327 }  )+$signed( -{ 2'b0,x328 }<<<3'd1 )+$signed( { 3'b0,x329 }<<<3'd2 )+$signed( { 3'b0,x331 }<<<3'd2 )+$signed( -{ 1'b0,x332 } )+$signed( { 3'b0,x333 }<<<3'd2 )+$signed( { 2'b0,x334 } <<<3'd1 )+$signed( -{ 3'b0,x335 }<<<3'd2)+$signed( -{ 3'b0,x336 }<<<3'd2)+$signed( -{ 1'b0,x337 } )+$signed( -{ 4'b0, x338 }<<<3'd3 )+$signed( { 2'b0,x339 } <<<3'd1 )+$signed( -{ 2'b0,x340 }<<<3'd1 )+$signed( -{ 2'b0,x342 }<<<3'd1 )+$signed( { 1'b0,x345 }  )+$signed( -{ 2'b0,x346 }<<<3'd1 )+$signed( { 3'b0,x347 }<<<3'd2 )+$signed( { 2'b0,x349 } <<<3'd1 )+$signed( -{ 5'b0,x351 }<<<3'd4 )+$signed( -{ 2'b0,x352 }<<<3'd1 )+$signed( -{ 2'b0,x353 }<<<3'd1 )+$signed( { 3'b0,x354 }<<<3'd2 )+$signed( { 2'b0,x355 } <<<3'd1 )+$signed( { 3'b0,x356 }<<<3'd2 )+$signed( { 3'b0,x357 }<<<3'd2 )+$signed( { 2'b0,x358 } <<<3'd1 )+$signed( -{ 1'b0,x359 } )+$signed( { 3'b0,x360 }<<<3'd2 )+$signed( { 1'b0,x361 }  )+$signed( { 2'b0,x363 } <<<3'd1 )+$signed( -{ 2'b0,x364 }<<<3'd1 )+$signed( -{ 3'b0,x365 }<<<3'd2)+$signed( -{ 2'b0,x366 }<<<3'd1 )+$signed( -{ 2'b0,x368 }<<<3'd1 )+$signed( { 1'b0,x369 }  )+$signed( { 4'b0,x370 }<<<3'd3 )+$signed( { 3'b0,x371 }<<<3'd2 )+$signed( -{ 1'b0,x372 } )+$signed( { 2'b0,x373 } <<<3'd1 )+$signed( { 1'b0,x374 }  )+$signed( -{ 3'b0,x375 }<<<3'd2)+$signed( -{ 3'b0,x376 }<<<3'd2)+$signed( -{ 2'b0,x377 }<<<3'd1 )+$signed( { 3'b0,x378 }<<<3'd2 )+$signed( { 1'b0,x379 }  )+$signed( -{ 1'b0,x381 } )+$signed( { 4'b0,x382 }<<<3'd3 )+$signed( { 4'b0,x383 }<<<3'd3 )+$signed( -{ 1'b0,x384 } )+$signed( { 3'b0,x385 }<<<3'd2 )+$signed( { 3'b0,x386 }<<<3'd2 )+$signed( { 2'b0,x387 } <<<3'd1 )+$signed( -{ 3'b0,x388 }<<<3'd2)+$signed( -{ 2'b0,x389 }<<<3'd1 )+$signed( -{ 4'b0, x390 }<<<3'd3 )+$signed( { 2'b0,x391 } <<<3'd1 )+$signed( { 3'b0,x392 }<<<3'd2 )+$signed( { 2'b0,x393 } <<<3'd1 )+$signed( { 1'b0,x394 }  )+$signed( { 3'b0,x395 }<<<3'd2 )+$signed( { 2'b0,x396 } <<<3'd1 )+$signed( -{ 2'b0,x398 }<<<3'd1 )+$signed( { 3'b0,x399 }<<<3'd2 )+$signed( -{ 3'b0,x400 }<<<3'd2)+$signed( -{ 2'b0,x402 }<<<3'd1 )+$signed( -{ 2'b0,x403 }<<<3'd1 )+$signed( -{ 1'b0,x404 } )+$signed( -{ 3'b0,x405 }<<<3'd2)+$signed( { 2'b0,x408 } <<<3'd1 )+$signed( { 1'b0,x409 }  )+$signed( { 3'b0,x410 }<<<3'd2 )+$signed( { 3'b0,x411 }<<<3'd2 )+$signed( { 3'b0,x412 }<<<3'd2 )+$signed( -{ 3'b0,x414 }<<<3'd2)+$signed( { 3'b0,x415 }<<<3'd2 )+$signed( { 3'b0,x416 }<<<3'd2 )+$signed( { 1'b0,x417 }  )+$signed( { 2'b0,x418 } <<<3'd1 )+$signed( -{ 2'b0,x419 }<<<3'd1 )+$signed( -{ 1'b0,x420 } )+$signed( { 2'b0,x421 } <<<3'd1 )+$signed( -{ 2'b0,x422 }<<<3'd1 )+$signed( { 3'b0,x423 }<<<3'd2 )+$signed( -{ 2'b0,x424 }<<<3'd1 )+$signed( -{ 1'b0,x425 } )+$signed( -{ 4'b0, x426 }<<<3'd3 )+$signed( { 3'b0,x427 }<<<3'd2 )+$signed( { 3'b0,x429 }<<<3'd2 )+$signed( -{ 3'b0,x430 }<<<3'd2)+$signed( -{ 3'b0,x433 }<<<3'd2)+$signed( -{ 1'b0,x434 } )+$signed( -{ 3'b0,x435 }<<<3'd2)+$signed( { 3'b0,x436 }<<<3'd2 )+$signed( { 3'b0,x437 }<<<3'd2 )+$signed( { 2'b0,x438 } <<<3'd1 )+$signed( -{ 3'b0,x439 }<<<3'd2)+$signed( { 2'b0,x441 } <<<3'd1 )+$signed( -{ 1'b0,x442 } )+$signed( { 3'b0,x443 }<<<3'd2 )+$signed( { 2'b0,x444 } <<<3'd1 )+$signed( -{ 1'b0,x445 } )+$signed( { 3'b0,x447 }<<<3'd2 )+$signed( -{ 2'b0,x448 }<<<3'd1 )+$signed( { 3'b0,x449 }<<<3'd2 )+$signed( { 1'b0,x450 }  )+$signed( -{ 1'b0,x451 } )+$signed( { 1'b0,x452 }  )+$signed( { 3'b0,x455 }<<<3'd2 )+$signed( -{ 2'b0,x456 }<<<3'd1 )+$signed( { 3'b0,x457 }<<<3'd2 )+$signed( { 2'b0,x458 } <<<3'd1 )+$signed( -{ 2'b0,x459 }<<<3'd1 )+$signed( { 2'b0,x460 } <<<3'd1 )+$signed( -{ 2'b0,x461 }<<<3'd1 )+$signed( { 2'b0,x462 } <<<3'd1 )+$signed( { 3'b0,x463 }<<<3'd2 )+$signed( -{ 1'b0,x465 } )+$signed( { 2'b0,x466 } <<<3'd1 )+$signed( -{ 1'b0,x467 } )+$signed( -{ 3'b0,x468 }<<<3'd2)+$signed( -{ 3'b0,x469 }<<<3'd2)+$signed( { 3'b0,x470 }<<<3'd2 )+$signed( -{ 2'b0,x471 }<<<3'd1 )+$signed( -{ 2'b0,x472 }<<<3'd1 )+$signed( -{ 2'b0,x473 }<<<3'd1 )+$signed( -{ 2'b0,x474 }<<<3'd1 )+$signed( { 2'b0,x475 } <<<3'd1 )+$signed( -{ 1'b0,x476 } )+$signed( -{ 2'b0,x477 }<<<3'd1 )+$signed( -{ 1'b0,x478 } )+$signed( -{ 3'b0,x480 }<<<3'd2)+$signed( -{ 1'b0,x481 } )+$signed( -{ 2'b0,x482 }<<<3'd1 )+$signed( { 3'b0,x483 }<<<3'd2 )+$signed( -{ 2'b0,x484 }<<<3'd1 )+$signed( { 2'b0,x485 } <<<3'd1 )+$signed( -{ 3'b0,x486 }<<<3'd2)+$signed( -{ 3'b0,x487 }<<<3'd2)+$signed( { 1'b0,x488 }  )+$signed( -{ 1'b0,x489 } )+$signed( -{ 1'b0,x490 } )+$signed( -{ 2'b0,x491 }<<<3'd1 )+$signed( { 3'b0,x492 }<<<3'd2 )+$signed( { 3'b0,x493 }<<<3'd2 )+$signed( -{ 2'b0,x494 }<<<3'd1 )+$signed( -{ 3'b0,x495 }<<<3'd2)+$signed(13'd8);
assign y1=temp_y[1][13] ==1'b1 ? 6'd0 :  
    temp_y[1][10] ==1'b1 ? 6'd63 : 
    temp_y[1][3]==1'b1 ? temp_y[1][9:4]+1'b1 : temp_y[1][9:4];
assign temp_y[2] = 
+$signed( -{ 2'b0,x0 }<<<3'd1 )+$signed( { 2'b0,x1 } <<<3'd1 )+$signed( -{ 2'b0,x3 }<<<3'd1 )+$signed( -{ 2'b0,x5 }<<<3'd1 )+$signed( { 3'b0,x7 }<<<3'd2 )+$signed( { 2'b0,x8 } <<<3'd1 )+$signed( -{ 2'b0,x10 }<<<3'd1 )+$signed( -{ 1'b0,x11 } )+$signed( -{ 2'b0,x12 }<<<3'd1 )+$signed( -{ 3'b0,x13 }<<<3'd2)+$signed( -{ 2'b0,x14 }<<<3'd1 )+$signed( { 2'b0,x16 } <<<3'd1 )+$signed( -{ 2'b0,x17 }<<<3'd1 )+$signed( { 2'b0,x18 } <<<3'd1 )+$signed( { 2'b0,x19 } <<<3'd1 )+$signed( -{ 1'b0,x20 } )+$signed( -{ 2'b0,x21 }<<<3'd1 )+$signed( { 2'b0,x22 } <<<3'd1 )+$signed( { 3'b0,x24 }<<<3'd2 )+$signed( { 2'b0,x25 } <<<3'd1 )+$signed( -{ 2'b0,x26 }<<<3'd1 )+$signed( -{ 2'b0,x27 }<<<3'd1 )+$signed( -{ 3'b0,x28 }<<<3'd2)+$signed( -{ 1'b0,x29 } )+$signed( -{ 3'b0,x30 }<<<3'd2)+$signed( -{ 1'b0,x31 } )+$signed( { 1'b0,x34 }  )+$signed( -{ 1'b0,x35 } )+$signed( -{ 3'b0,x36 }<<<3'd2)+$signed( { 1'b0,x39 }  )+$signed( { 1'b0,x40 }  )+$signed( -{ 1'b0,x41 } )+$signed( -{ 1'b0,x42 } )+$signed( { 3'b0,x43 }<<<3'd2 )+$signed( -{ 3'b0,x45 }<<<3'd2)+$signed( { 2'b0,x46 } <<<3'd1 )+$signed( -{ 2'b0,x47 }<<<3'd1 )+$signed( -{ 2'b0,x48 }<<<3'd1 )+$signed( -{ 2'b0,x49 }<<<3'd1 )+$signed( { 3'b0,x50 }<<<3'd2 )+$signed( { 2'b0,x51 } <<<3'd1 )+$signed( { 3'b0,x53 }<<<3'd2 )+$signed( -{ 2'b0,x54 }<<<3'd1 )+$signed( { 2'b0,x55 } <<<3'd1 )+$signed( -{ 2'b0,x58 }<<<3'd1 )+$signed( -{ 1'b0,x59 } )+$signed( { 2'b0,x60 } <<<3'd1 )+$signed( { 3'b0,x61 }<<<3'd2 )+$signed( { 1'b0,x62 }  )+$signed( -{ 1'b0,x63 } )+$signed( { 2'b0,x64 } <<<3'd1 )+$signed( -{ 2'b0,x65 }<<<3'd1 )+$signed( { 3'b0,x66 }<<<3'd2 )+$signed( -{ 2'b0,x67 }<<<3'd1 )+$signed( -{ 2'b0,x70 }<<<3'd1 )+$signed( -{ 1'b0,x71 } )+$signed( -{ 4'b0, x72 }<<<3'd3 )+$signed( { 2'b0,x73 } <<<3'd1 )+$signed( { 1'b0,x74 }  )+$signed( { 3'b0,x75 }<<<3'd2 )+$signed( { 1'b0,x77 }  )+$signed( -{ 2'b0,x79 }<<<3'd1 )+$signed( { 2'b0,x80 } <<<3'd1 )+$signed( { 2'b0,x81 } <<<3'd1 )+$signed( { 3'b0,x82 }<<<3'd2 )+$signed( -{ 1'b0,x83 } )+$signed( -{ 3'b0,x84 }<<<3'd2)+$signed( -{ 3'b0,x85 }<<<3'd2)+$signed( -{ 1'b0,x86 } )+$signed( { 1'b0,x87 }  )+$signed( { 1'b0,x88 }  )+$signed( -{ 3'b0,x90 }<<<3'd2)+$signed( { 3'b0,x91 }<<<3'd2 )+$signed( { 3'b0,x92 }<<<3'd2 )+$signed( { 3'b0,x93 }<<<3'd2 )+$signed( { 3'b0,x94 }<<<3'd2 )+$signed( -{ 2'b0,x95 }<<<3'd1 )+$signed( -{ 2'b0,x96 }<<<3'd1 )+$signed( { 3'b0,x97 }<<<3'd2 )+$signed( { 1'b0,x98 }  )+$signed( { 1'b0,x99 }  )+$signed( -{ 2'b0,x100 }<<<3'd1 )+$signed( -{ 2'b0,x101 }<<<3'd1 )+$signed( { 3'b0,x102 }<<<3'd2 )+$signed( { 1'b0,x103 }  )+$signed( -{ 2'b0,x104 }<<<3'd1 )+$signed( { 2'b0,x106 } <<<3'd1 )+$signed( -{ 2'b0,x108 }<<<3'd1 )+$signed( { 3'b0,x109 }<<<3'd2 )+$signed( { 2'b0,x110 } <<<3'd1 )+$signed( -{ 3'b0,x111 }<<<3'd2)+$signed( -{ 2'b0,x113 }<<<3'd1 )+$signed( -{ 3'b0,x114 }<<<3'd2)+$signed( { 4'b0,x115 }<<<3'd3 )+$signed( { 2'b0,x116 } <<<3'd1 )+$signed( -{ 2'b0,x117 }<<<3'd1 )+$signed( -{ 2'b0,x118 }<<<3'd1 )+$signed( { 1'b0,x119 }  )+$signed( { 2'b0,x120 } <<<3'd1 )+$signed( { 2'b0,x121 } <<<3'd1 )+$signed( -{ 3'b0,x122 }<<<3'd2)+$signed( { 3'b0,x123 }<<<3'd2 )+$signed( -{ 1'b0,x124 } )+$signed( -{ 1'b0,x125 } )+$signed( -{ 1'b0,x126 } )+$signed( { 2'b0,x129 } <<<3'd1 )+$signed( { 1'b0,x130 }  )+$signed( { 3'b0,x131 }<<<3'd2 )+$signed( { 1'b0,x132 }  )+$signed( { 3'b0,x133 }<<<3'd2 )+$signed( { 1'b0,x134 }  )+$signed( { 1'b0,x135 }  )+$signed( { 3'b0,x136 }<<<3'd2 )+$signed( { 2'b0,x137 } <<<3'd1 )+$signed( -{ 3'b0,x138 }<<<3'd2)+$signed( -{ 3'b0,x139 }<<<3'd2)+$signed( { 1'b0,x141 }  )+$signed( -{ 2'b0,x142 }<<<3'd1 )+$signed( { 1'b0,x143 }  )+$signed( { 1'b0,x144 }  )+$signed( { 2'b0,x145 } <<<3'd1 )+$signed( { 1'b0,x147 }  )+$signed( -{ 2'b0,x148 }<<<3'd1 )+$signed( -{ 1'b0,x149 } )+$signed( -{ 2'b0,x151 }<<<3'd1 )+$signed( { 3'b0,x152 }<<<3'd2 )+$signed( -{ 2'b0,x153 }<<<3'd1 )+$signed( { 3'b0,x154 }<<<3'd2 )+$signed( { 1'b0,x156 }  )+$signed( -{ 2'b0,x157 }<<<3'd1 )+$signed( -{ 2'b0,x158 }<<<3'd1 )+$signed( -{ 2'b0,x159 }<<<3'd1 )+$signed( -{ 2'b0,x160 }<<<3'd1 )+$signed( { 2'b0,x161 } <<<3'd1 )+$signed( { 2'b0,x162 } <<<3'd1 )+$signed( { 3'b0,x164 }<<<3'd2 )+$signed( { 2'b0,x165 } <<<3'd1 )+$signed( { 1'b0,x166 }  )+$signed( { 2'b0,x167 } <<<3'd1 )+$signed( -{ 2'b0,x168 }<<<3'd1 )+$signed( -{ 1'b0,x169 } )+$signed( -{ 1'b0,x170 } )+$signed( -{ 2'b0,x171 }<<<3'd1 )+$signed( { 3'b0,x172 }<<<3'd2 )+$signed( { 2'b0,x173 } <<<3'd1 )+$signed( -{ 2'b0,x174 }<<<3'd1 )+$signed( -{ 1'b0,x175 } )+$signed( -{ 1'b0,x176 } )+$signed( { 1'b0,x177 }  )+$signed( -{ 2'b0,x178 }<<<3'd1 )+$signed( { 3'b0,x179 }<<<3'd2 )+$signed( { 1'b0,x180 }  )+$signed( { 2'b0,x181 } <<<3'd1 )+$signed( { 2'b0,x182 } <<<3'd1 )+$signed( { 1'b0,x183 }  )+$signed( { 1'b0,x184 }  )+$signed( { 2'b0,x185 } <<<3'd1 )+$signed( -{ 1'b0,x186 } )+$signed( { 3'b0,x187 }<<<3'd2 )+$signed( -{ 2'b0,x188 }<<<3'd1 )+$signed( -{ 3'b0,x190 }<<<3'd2)+$signed( { 2'b0,x191 } <<<3'd1 )+$signed( -{ 3'b0,x192 }<<<3'd2)+$signed( -{ 2'b0,x193 }<<<3'd1 )+$signed( -{ 1'b0,x194 } )+$signed( { 3'b0,x195 }<<<3'd2 )+$signed( -{ 2'b0,x196 }<<<3'd1 )+$signed( { 3'b0,x197 }<<<3'd2 )+$signed( { 2'b0,x198 } <<<3'd1 )+$signed( { 2'b0,x199 } <<<3'd1 )+$signed( -{ 2'b0,x200 }<<<3'd1 )+$signed( { 3'b0,x201 }<<<3'd2 )+$signed( -{ 3'b0,x205 }<<<3'd2)+$signed( { 2'b0,x206 } <<<3'd1 )+$signed( { 2'b0,x208 } <<<3'd1 )+$signed( { 2'b0,x210 } <<<3'd1 )+$signed( -{ 2'b0,x211 }<<<3'd1 )+$signed( { 1'b0,x212 }  )+$signed( { 2'b0,x213 } <<<3'd1 )+$signed( -{ 2'b0,x214 }<<<3'd1 )+$signed( { 3'b0,x215 }<<<3'd2 )+$signed( { 3'b0,x216 }<<<3'd2 )+$signed( { 3'b0,x217 }<<<3'd2 )+$signed( { 3'b0,x218 }<<<3'd2 )+$signed( -{ 3'b0,x219 }<<<3'd2)+$signed( -{ 3'b0,x220 }<<<3'd2)+$signed( { 1'b0,x221 }  )+$signed( { 3'b0,x222 }<<<3'd2 )+$signed( -{ 2'b0,x223 }<<<3'd1 )+$signed( { 3'b0,x224 }<<<3'd2 )+$signed( { 2'b0,x226 } <<<3'd1 )+$signed( -{ 1'b0,x227 } )+$signed( -{ 1'b0,x228 } )+$signed( { 3'b0,x229 }<<<3'd2 )+$signed( -{ 1'b0,x230 } )+$signed( -{ 3'b0,x231 }<<<3'd2)+$signed( { 1'b0,x232 }  )+$signed( -{ 1'b0,x233 } )+$signed( { 3'b0,x235 }<<<3'd2 )+$signed( { 4'b0,x236 }<<<3'd3 )+$signed( -{ 2'b0,x237 }<<<3'd1 )+$signed( { 2'b0,x238 } <<<3'd1 )+$signed( { 1'b0,x240 }  )+$signed( -{ 3'b0,x241 }<<<3'd2)+$signed( { 1'b0,x242 }  )+$signed( -{ 2'b0,x243 }<<<3'd1 )+$signed( { 1'b0,x244 }  )+$signed( -{ 1'b0,x245 } )+$signed( -{ 2'b0,x246 }<<<3'd1 )+$signed( -{ 3'b0,x247 }<<<3'd2)+$signed( -{ 3'b0,x248 }<<<3'd2)+$signed( { 3'b0,x249 }<<<3'd2 )+$signed( -{ 3'b0,x250 }<<<3'd2)+$signed( { 2'b0,x251 } <<<3'd1 )+$signed( -{ 2'b0,x252 }<<<3'd1 )+$signed( { 1'b0,x253 }  )+$signed( { 4'b0,x254 }<<<3'd3 )+$signed( { 2'b0,x255 } <<<3'd1 )+$signed( { 2'b0,x256 } <<<3'd1 )+$signed( -{ 1'b0,x257 } )+$signed( { 1'b0,x258 }  )+$signed( -{ 2'b0,x259 }<<<3'd1 )+$signed( { 2'b0,x260 } <<<3'd1 )+$signed( -{ 3'b0,x261 }<<<3'd2)+$signed( -{ 2'b0,x262 }<<<3'd1 )+$signed( -{ 2'b0,x264 }<<<3'd1 )+$signed( -{ 3'b0,x265 }<<<3'd2)+$signed( -{ 1'b0,x266 } )+$signed( { 3'b0,x267 }<<<3'd2 )+$signed( -{ 2'b0,x268 }<<<3'd1 )+$signed( { 2'b0,x269 } <<<3'd1 )+$signed( -{ 1'b0,x272 } )+$signed( { 2'b0,x273 } <<<3'd1 )+$signed( -{ 3'b0,x274 }<<<3'd2)+$signed( { 2'b0,x275 } <<<3'd1 )+$signed( { 3'b0,x276 }<<<3'd2 )+$signed( -{ 3'b0,x277 }<<<3'd2)+$signed( { 3'b0,x278 }<<<3'd2 )+$signed( { 2'b0,x280 } <<<3'd1 )+$signed( -{ 3'b0,x281 }<<<3'd2)+$signed( { 1'b0,x282 }  )+$signed( -{ 1'b0,x283 } )+$signed( { 2'b0,x284 } <<<3'd1 )+$signed( -{ 1'b0,x286 } )+$signed( { 3'b0,x288 }<<<3'd2 )+$signed( { 3'b0,x289 }<<<3'd2 )+$signed( { 2'b0,x290 } <<<3'd1 )+$signed( -{ 1'b0,x291 } )+$signed( -{ 2'b0,x292 }<<<3'd1 )+$signed( -{ 2'b0,x293 }<<<3'd1 )+$signed( -{ 2'b0,x294 }<<<3'd1 )+$signed( { 3'b0,x296 }<<<3'd2 )+$signed( -{ 3'b0,x297 }<<<3'd2)+$signed( -{ 1'b0,x298 } )+$signed( -{ 3'b0,x299 }<<<3'd2)+$signed( -{ 1'b0,x300 } )+$signed( { 3'b0,x301 }<<<3'd2 )+$signed( { 2'b0,x302 } <<<3'd1 )+$signed( -{ 2'b0,x303 }<<<3'd1 )+$signed( -{ 2'b0,x304 }<<<3'd1 )+$signed( -{ 2'b0,x305 }<<<3'd1 )+$signed( -{ 2'b0,x306 }<<<3'd1 )+$signed( { 1'b0,x308 }  )+$signed( -{ 1'b0,x309 } )+$signed( -{ 1'b0,x310 } )+$signed( { 2'b0,x312 } <<<3'd1 )+$signed( { 2'b0,x313 } <<<3'd1 )+$signed( -{ 2'b0,x314 }<<<3'd1 )+$signed( { 1'b0,x315 }  )+$signed( { 1'b0,x316 }  )+$signed( { 3'b0,x317 }<<<3'd2 )+$signed( { 1'b0,x318 }  )+$signed( -{ 3'b0,x319 }<<<3'd2)+$signed( { 2'b0,x320 } <<<3'd1 )+$signed( -{ 1'b0,x321 } )+$signed( -{ 3'b0,x322 }<<<3'd2)+$signed( -{ 1'b0,x323 } )+$signed( -{ 3'b0,x325 }<<<3'd2)+$signed( { 1'b0,x326 }  )+$signed( { 3'b0,x327 }<<<3'd2 )+$signed( -{ 1'b0,x328 } )+$signed( -{ 2'b0,x329 }<<<3'd1 )+$signed( { 2'b0,x330 } <<<3'd1 )+$signed( { 4'b0,x331 }<<<3'd3 )+$signed( -{ 3'b0,x332 }<<<3'd2)+$signed( { 1'b0,x333 }  )+$signed( -{ 2'b0,x334 }<<<3'd1 )+$signed( { 2'b0,x335 } <<<3'd1 )+$signed( { 1'b0,x336 }  )+$signed( { 2'b0,x337 } <<<3'd1 )+$signed( -{ 2'b0,x339 }<<<3'd1 )+$signed( -{ 3'b0,x341 }<<<3'd2)+$signed( -{ 1'b0,x342 } )+$signed( { 2'b0,x343 } <<<3'd1 )+$signed( -{ 1'b0,x344 } )+$signed( -{ 3'b0,x345 }<<<3'd2)+$signed( { 1'b0,x346 }  )+$signed( -{ 3'b0,x347 }<<<3'd2)+$signed( { 2'b0,x348 } <<<3'd1 )+$signed( { 1'b0,x350 }  )+$signed( { 1'b0,x352 }  )+$signed( -{ 3'b0,x353 }<<<3'd2)+$signed( { 2'b0,x354 } <<<3'd1 )+$signed( { 3'b0,x355 }<<<3'd2 )+$signed( { 3'b0,x356 }<<<3'd2 )+$signed( { 3'b0,x357 }<<<3'd2 )+$signed( { 3'b0,x358 }<<<3'd2 )+$signed( { 3'b0,x359 }<<<3'd2 )+$signed( { 2'b0,x360 } <<<3'd1 )+$signed( { 4'b0,x361 }<<<3'd3 )+$signed( { 2'b0,x362 } <<<3'd1 )+$signed( -{ 1'b0,x363 } )+$signed( { 3'b0,x364 }<<<3'd2 )+$signed( { 3'b0,x365 }<<<3'd2 )+$signed( { 1'b0,x366 }  )+$signed( -{ 1'b0,x367 } )+$signed( { 1'b0,x368 }  )+$signed( { 2'b0,x370 } <<<3'd1 )+$signed( { 3'b0,x371 }<<<3'd2 )+$signed( { 2'b0,x372 } <<<3'd1 )+$signed( -{ 1'b0,x373 } )+$signed( { 2'b0,x374 } <<<3'd1 )+$signed( { 2'b0,x375 } <<<3'd1 )+$signed( { 2'b0,x376 } <<<3'd1 )+$signed( { 2'b0,x377 } <<<3'd1 )+$signed( { 3'b0,x378 }<<<3'd2 )+$signed( { 1'b0,x379 }  )+$signed( -{ 3'b0,x380 }<<<3'd2)+$signed( { 2'b0,x381 } <<<3'd1 )+$signed( -{ 1'b0,x382 } )+$signed( -{ 3'b0,x384 }<<<3'd2)+$signed( { 2'b0,x385 } <<<3'd1 )+$signed( -{ 3'b0,x386 }<<<3'd2)+$signed( { 2'b0,x388 } <<<3'd1 )+$signed( { 2'b0,x389 } <<<3'd1 )+$signed( -{ 2'b0,x390 }<<<3'd1 )+$signed( { 3'b0,x391 }<<<3'd2 )+$signed( { 2'b0,x392 } <<<3'd1 )+$signed( -{ 3'b0,x393 }<<<3'd2)+$signed( { 3'b0,x394 }<<<3'd2 )+$signed( { 1'b0,x395 }  )+$signed( { 1'b0,x396 }  )+$signed( -{ 3'b0,x397 }<<<3'd2)+$signed( -{ 1'b0,x398 } )+$signed( -{ 3'b0,x399 }<<<3'd2)+$signed( -{ 2'b0,x400 }<<<3'd1 )+$signed( { 4'b0,x403 }<<<3'd3 )+$signed( -{ 3'b0,x404 }<<<3'd2)+$signed( -{ 2'b0,x405 }<<<3'd1 )+$signed( { 3'b0,x406 }<<<3'd2 )+$signed( { 3'b0,x407 }<<<3'd2 )+$signed( { 4'b0,x408 }<<<3'd3 )+$signed( { 1'b0,x409 }  )+$signed( { 3'b0,x411 }<<<3'd2 )+$signed( { 2'b0,x412 } <<<3'd1 )+$signed( { 1'b0,x413 }  )+$signed( -{ 1'b0,x414 } )+$signed( -{ 1'b0,x415 } )+$signed( { 3'b0,x416 }<<<3'd2 )+$signed( -{ 2'b0,x417 }<<<3'd1 )+$signed( { 3'b0,x418 }<<<3'd2 )+$signed( { 2'b0,x419 } <<<3'd1 )+$signed( { 3'b0,x420 }<<<3'd2 )+$signed( { 2'b0,x421 } <<<3'd1 )+$signed( { 2'b0,x422 } <<<3'd1 )+$signed( -{ 2'b0,x423 }<<<3'd1 )+$signed( -{ 1'b0,x424 } )+$signed( -{ 2'b0,x425 }<<<3'd1 )+$signed( { 3'b0,x426 }<<<3'd2 )+$signed( { 2'b0,x428 } <<<3'd1 )+$signed( -{ 2'b0,x429 }<<<3'd1 )+$signed( { 2'b0,x430 } <<<3'd1 )+$signed( -{ 1'b0,x431 } )+$signed( { 2'b0,x432 } <<<3'd1 )+$signed( { 4'b0,x433 }<<<3'd3 )+$signed( -{ 1'b0,x434 } )+$signed( { 1'b0,x435 }  )+$signed( -{ 1'b0,x436 } )+$signed( -{ 2'b0,x437 }<<<3'd1 )+$signed( -{ 2'b0,x438 }<<<3'd1 )+$signed( -{ 2'b0,x439 }<<<3'd1 )+$signed( { 2'b0,x440 } <<<3'd1 )+$signed( { 1'b0,x441 }  )+$signed( -{ 3'b0,x442 }<<<3'd2)+$signed( { 2'b0,x443 } <<<3'd1 )+$signed( { 4'b0,x444 }<<<3'd3 )+$signed( -{ 2'b0,x445 }<<<3'd1 )+$signed( -{ 3'b0,x447 }<<<3'd2)+$signed( -{ 2'b0,x448 }<<<3'd1 )+$signed( -{ 1'b0,x449 } )+$signed( { 1'b0,x450 }  )+$signed( -{ 2'b0,x451 }<<<3'd1 )+$signed( -{ 2'b0,x452 }<<<3'd1 )+$signed( -{ 1'b0,x453 } )+$signed( { 2'b0,x455 } <<<3'd1 )+$signed( -{ 2'b0,x456 }<<<3'd1 )+$signed( -{ 1'b0,x457 } )+$signed( -{ 1'b0,x458 } )+$signed( { 4'b0,x459 }<<<3'd3 )+$signed( -{ 1'b0,x460 } )+$signed( -{ 2'b0,x462 }<<<3'd1 )+$signed( { 3'b0,x463 }<<<3'd2 )+$signed( -{ 2'b0,x464 }<<<3'd1 )+$signed( { 1'b0,x465 }  )+$signed( { 3'b0,x467 }<<<3'd2 )+$signed( { 2'b0,x468 } <<<3'd1 )+$signed( -{ 2'b0,x469 }<<<3'd1 )+$signed( -{ 3'b0,x470 }<<<3'd2)+$signed( { 3'b0,x472 }<<<3'd2 )+$signed( -{ 1'b0,x473 } )+$signed( { 2'b0,x474 } <<<3'd1 )+$signed( -{ 3'b0,x475 }<<<3'd2)+$signed( { 3'b0,x476 }<<<3'd2 )+$signed( -{ 1'b0,x477 } )+$signed( { 1'b0,x478 }  )+$signed( { 2'b0,x479 } <<<3'd1 )+$signed( { 4'b0,x480 }<<<3'd3 )+$signed( -{ 2'b0,x481 }<<<3'd1 )+$signed( -{ 2'b0,x482 }<<<3'd1 )+$signed( -{ 3'b0,x483 }<<<3'd2)+$signed( -{ 2'b0,x484 }<<<3'd1 )+$signed( { 1'b0,x485 }  )+$signed( { 1'b0,x486 }  )+$signed( { 3'b0,x487 }<<<3'd2 )+$signed( -{ 1'b0,x488 } )+$signed( -{ 1'b0,x490 } )+$signed( { 2'b0,x492 } <<<3'd1 )+$signed( { 3'b0,x493 }<<<3'd2 )+$signed( { 1'b0,x495 }  )+$signed(13'd32);
assign y2=temp_y[2][13] ==1'b1 ? 6'd0 :  
    temp_y[2][10] ==1'b1 ? 6'd63 : 
    temp_y[2][3]==1'b1 ? temp_y[2][9:4]+1'b1 : temp_y[2][9:4];
assign temp_y[3] = 
+$signed( -{ 1'b0,x0 } )+$signed( { 2'b0,x1 } <<<3'd1 )+$signed( { 1'b0,x2 }  )+$signed( { 4'b0,x3 }<<<3'd3 )+$signed( { 2'b0,x4 } <<<3'd1 )+$signed( -{ 3'b0,x5 }<<<3'd2)+$signed( { 1'b0,x6 }  )+$signed( -{ 3'b0,x7 }<<<3'd2)+$signed( { 1'b0,x8 }  )+$signed( -{ 2'b0,x9 }<<<3'd1 )+$signed( { 1'b0,x10 }  )+$signed( -{ 3'b0,x12 }<<<3'd2)+$signed( -{ 1'b0,x13 } )+$signed( -{ 2'b0,x14 }<<<3'd1 )+$signed( { 3'b0,x16 }<<<3'd2 )+$signed( { 2'b0,x17 } <<<3'd1 )+$signed( { 3'b0,x18 }<<<3'd2 )+$signed( -{ 1'b0,x19 } )+$signed( -{ 2'b0,x20 }<<<3'd1 )+$signed( { 2'b0,x21 } <<<3'd1 )+$signed( { 3'b0,x22 }<<<3'd2 )+$signed( -{ 1'b0,x24 } )+$signed( -{ 2'b0,x25 }<<<3'd1 )+$signed( -{ 1'b0,x26 } )+$signed( -{ 2'b0,x27 }<<<3'd1 )+$signed( -{ 3'b0,x28 }<<<3'd2)+$signed( { 1'b0,x29 }  )+$signed( { 3'b0,x30 }<<<3'd2 )+$signed( { 2'b0,x31 } <<<3'd1 )+$signed( { 1'b0,x32 }  )+$signed( -{ 3'b0,x33 }<<<3'd2)+$signed( -{ 1'b0,x34 } )+$signed( { 2'b0,x35 } <<<3'd1 )+$signed( -{ 1'b0,x36 } )+$signed( -{ 2'b0,x37 }<<<3'd1 )+$signed( -{ 3'b0,x38 }<<<3'd2)+$signed( { 3'b0,x39 }<<<3'd2 )+$signed( { 3'b0,x40 }<<<3'd2 )+$signed( { 1'b0,x41 }  )+$signed( { 1'b0,x42 }  )+$signed( { 1'b0,x44 }  )+$signed( -{ 3'b0,x45 }<<<3'd2)+$signed( -{ 3'b0,x46 }<<<3'd2)+$signed( { 2'b0,x47 } <<<3'd1 )+$signed( { 2'b0,x49 } <<<3'd1 )+$signed( { 2'b0,x50 } <<<3'd1 )+$signed( -{ 3'b0,x51 }<<<3'd2)+$signed( { 1'b0,x52 }  )+$signed( { 2'b0,x53 } <<<3'd1 )+$signed( { 2'b0,x54 } <<<3'd1 )+$signed( { 2'b0,x55 } <<<3'd1 )+$signed( -{ 2'b0,x56 }<<<3'd1 )+$signed( { 3'b0,x57 }<<<3'd2 )+$signed( { 3'b0,x58 }<<<3'd2 )+$signed( -{ 2'b0,x61 }<<<3'd1 )+$signed( { 1'b0,x62 }  )+$signed( { 2'b0,x63 } <<<3'd1 )+$signed( { 3'b0,x64 }<<<3'd2 )+$signed( { 2'b0,x65 } <<<3'd1 )+$signed( { 1'b0,x67 }  )+$signed( { 2'b0,x68 } <<<3'd1 )+$signed( -{ 3'b0,x69 }<<<3'd2)+$signed( { 3'b0,x70 }<<<3'd2 )+$signed( { 2'b0,x71 } <<<3'd1 )+$signed( -{ 2'b0,x72 }<<<3'd1 )+$signed( -{ 2'b0,x73 }<<<3'd1 )+$signed( { 2'b0,x74 } <<<3'd1 )+$signed( { 3'b0,x75 }<<<3'd2 )+$signed( { 3'b0,x76 }<<<3'd2 )+$signed( -{ 2'b0,x77 }<<<3'd1 )+$signed( { 1'b0,x79 }  )+$signed( -{ 1'b0,x80 } )+$signed( -{ 2'b0,x81 }<<<3'd1 )+$signed( -{ 1'b0,x82 } )+$signed( -{ 2'b0,x84 }<<<3'd1 )+$signed( -{ 2'b0,x85 }<<<3'd1 )+$signed( { 2'b0,x86 } <<<3'd1 )+$signed( { 2'b0,x87 } <<<3'd1 )+$signed( -{ 1'b0,x88 } )+$signed( -{ 2'b0,x89 }<<<3'd1 )+$signed( { 1'b0,x90 }  )+$signed( -{ 1'b0,x91 } )+$signed( { 3'b0,x92 }<<<3'd2 )+$signed( { 2'b0,x93 } <<<3'd1 )+$signed( { 4'b0,x94 }<<<3'd3 )+$signed( { 3'b0,x95 }<<<3'd2 )+$signed( -{ 2'b0,x96 }<<<3'd1 )+$signed( { 2'b0,x97 } <<<3'd1 )+$signed( -{ 3'b0,x98 }<<<3'd2)+$signed( -{ 2'b0,x99 }<<<3'd1 )+$signed( -{ 2'b0,x100 }<<<3'd1 )+$signed( { 2'b0,x101 } <<<3'd1 )+$signed( { 3'b0,x102 }<<<3'd2 )+$signed( { 2'b0,x103 } <<<3'd1 )+$signed( -{ 3'b0,x104 }<<<3'd2)+$signed( { 2'b0,x105 } <<<3'd1 )+$signed( { 2'b0,x106 } <<<3'd1 )+$signed( { 2'b0,x107 } <<<3'd1 )+$signed( -{ 1'b0,x108 } )+$signed( { 1'b0,x109 }  )+$signed( { 3'b0,x110 }<<<3'd2 )+$signed( { 2'b0,x111 } <<<3'd1 )+$signed( { 4'b0,x112 }<<<3'd3 )+$signed( { 3'b0,x113 }<<<3'd2 )+$signed( { 2'b0,x114 } <<<3'd1 )+$signed( -{ 1'b0,x115 } )+$signed( -{ 2'b0,x116 }<<<3'd1 )+$signed( -{ 2'b0,x117 }<<<3'd1 )+$signed( -{ 3'b0,x118 }<<<3'd2)+$signed( { 2'b0,x119 } <<<3'd1 )+$signed( { 2'b0,x120 } <<<3'd1 )+$signed( { 2'b0,x121 } <<<3'd1 )+$signed( -{ 1'b0,x122 } )+$signed( { 3'b0,x123 }<<<3'd2 )+$signed( { 1'b0,x124 }  )+$signed( { 1'b0,x125 }  )+$signed( { 2'b0,x126 } <<<3'd1 )+$signed( -{ 1'b0,x127 } )+$signed( { 1'b0,x128 }  )+$signed( { 3'b0,x129 }<<<3'd2 )+$signed( { 1'b0,x130 }  )+$signed( -{ 2'b0,x131 }<<<3'd1 )+$signed( -{ 2'b0,x133 }<<<3'd1 )+$signed( { 2'b0,x134 } <<<3'd1 )+$signed( { 1'b0,x135 }  )+$signed( { 2'b0,x136 } <<<3'd1 )+$signed( -{ 2'b0,x139 }<<<3'd1 )+$signed( -{ 2'b0,x140 }<<<3'd1 )+$signed( { 2'b0,x141 } <<<3'd1 )+$signed( { 2'b0,x142 } <<<3'd1 )+$signed( { 2'b0,x144 } <<<3'd1 )+$signed( -{ 2'b0,x145 }<<<3'd1 )+$signed( -{ 1'b0,x146 } )+$signed( { 2'b0,x147 } <<<3'd1 )+$signed( { 1'b0,x148 }  )+$signed( -{ 2'b0,x149 }<<<3'd1 )+$signed( -{ 2'b0,x150 }<<<3'd1 )+$signed( { 2'b0,x151 } <<<3'd1 )+$signed( -{ 1'b0,x152 } )+$signed( -{ 3'b0,x153 }<<<3'd2)+$signed( -{ 1'b0,x154 } )+$signed( { 2'b0,x155 } <<<3'd1 )+$signed( { 3'b0,x156 }<<<3'd2 )+$signed( -{ 2'b0,x157 }<<<3'd1 )+$signed( { 2'b0,x158 } <<<3'd1 )+$signed( -{ 2'b0,x160 }<<<3'd1 )+$signed( -{ 3'b0,x162 }<<<3'd2)+$signed( -{ 2'b0,x164 }<<<3'd1 )+$signed( { 3'b0,x165 }<<<3'd2 )+$signed( { 3'b0,x166 }<<<3'd2 )+$signed( -{ 1'b0,x167 } )+$signed( { 1'b0,x168 }  )+$signed( -{ 2'b0,x169 }<<<3'd1 )+$signed( { 1'b0,x170 }  )+$signed( { 2'b0,x172 } <<<3'd1 )+$signed( { 3'b0,x173 }<<<3'd2 )+$signed( { 3'b0,x174 }<<<3'd2 )+$signed( { 3'b0,x175 }<<<3'd2 )+$signed( { 3'b0,x176 }<<<3'd2 )+$signed( { 2'b0,x177 } <<<3'd1 )+$signed( { 2'b0,x178 } <<<3'd1 )+$signed( { 4'b0,x179 }<<<3'd3 )+$signed( -{ 1'b0,x181 } )+$signed( { 2'b0,x182 } <<<3'd1 )+$signed( { 2'b0,x183 } <<<3'd1 )+$signed( { 2'b0,x184 } <<<3'd1 )+$signed( -{ 1'b0,x185 } )+$signed( -{ 2'b0,x186 }<<<3'd1 )+$signed( -{ 3'b0,x187 }<<<3'd2)+$signed( -{ 2'b0,x188 }<<<3'd1 )+$signed( { 3'b0,x189 }<<<3'd2 )+$signed( { 3'b0,x191 }<<<3'd2 )+$signed( { 3'b0,x192 }<<<3'd2 )+$signed( { 3'b0,x193 }<<<3'd2 )+$signed( { 2'b0,x194 } <<<3'd1 )+$signed( -{ 1'b0,x195 } )+$signed( { 1'b0,x196 }  )+$signed( { 3'b0,x197 }<<<3'd2 )+$signed( -{ 1'b0,x198 } )+$signed( -{ 1'b0,x199 } )+$signed( -{ 2'b0,x200 }<<<3'd1 )+$signed( { 2'b0,x201 } <<<3'd1 )+$signed( -{ 2'b0,x203 }<<<3'd1 )+$signed( -{ 1'b0,x204 } )+$signed( -{ 2'b0,x205 }<<<3'd1 )+$signed( -{ 2'b0,x206 }<<<3'd1 )+$signed( -{ 2'b0,x207 }<<<3'd1 )+$signed( { 2'b0,x209 } <<<3'd1 )+$signed( { 3'b0,x210 }<<<3'd2 )+$signed( { 2'b0,x211 } <<<3'd1 )+$signed( { 3'b0,x212 }<<<3'd2 )+$signed( { 1'b0,x213 }  )+$signed( { 2'b0,x214 } <<<3'd1 )+$signed( { 3'b0,x215 }<<<3'd2 )+$signed( -{ 2'b0,x217 }<<<3'd1 )+$signed( { 2'b0,x219 } <<<3'd1 )+$signed( { 2'b0,x220 } <<<3'd1 )+$signed( -{ 3'b0,x221 }<<<3'd2)+$signed( { 2'b0,x222 } <<<3'd1 )+$signed( -{ 3'b0,x223 }<<<3'd2)+$signed( -{ 1'b0,x224 } )+$signed( -{ 1'b0,x225 } )+$signed( { 2'b0,x226 } <<<3'd1 )+$signed( { 1'b0,x227 }  )+$signed( { 1'b0,x228 }  )+$signed( { 1'b0,x229 }  )+$signed( { 1'b0,x230 }  )+$signed( { 2'b0,x231 } <<<3'd1 )+$signed( -{ 2'b0,x233 }<<<3'd1 )+$signed( -{ 1'b0,x234 } )+$signed( { 2'b0,x235 } <<<3'd1 )+$signed( -{ 2'b0,x236 }<<<3'd1 )+$signed( { 2'b0,x237 } <<<3'd1 )+$signed( { 3'b0,x238 }<<<3'd2 )+$signed( { 1'b0,x239 }  )+$signed( -{ 1'b0,x240 } )+$signed( -{ 2'b0,x242 }<<<3'd1 )+$signed( -{ 2'b0,x244 }<<<3'd1 )+$signed( -{ 1'b0,x246 } )+$signed( { 2'b0,x247 } <<<3'd1 )+$signed( -{ 1'b0,x248 } )+$signed( { 4'b0,x250 }<<<3'd3 )+$signed( -{ 2'b0,x251 }<<<3'd1 )+$signed( { 1'b0,x253 }  )+$signed( { 1'b0,x254 }  )+$signed( -{ 2'b0,x255 }<<<3'd1 )+$signed( { 2'b0,x256 } <<<3'd1 )+$signed( { 2'b0,x257 } <<<3'd1 )+$signed( -{ 1'b0,x259 } )+$signed( -{ 2'b0,x260 }<<<3'd1 )+$signed( -{ 1'b0,x261 } )+$signed( -{ 2'b0,x262 }<<<3'd1 )+$signed( { 1'b0,x266 }  )+$signed( -{ 2'b0,x267 }<<<3'd1 )+$signed( { 3'b0,x268 }<<<3'd2 )+$signed( { 2'b0,x269 } <<<3'd1 )+$signed( { 1'b0,x270 }  )+$signed( { 2'b0,x271 } <<<3'd1 )+$signed( -{ 2'b0,x272 }<<<3'd1 )+$signed( { 3'b0,x273 }<<<3'd2 )+$signed( { 2'b0,x274 } <<<3'd1 )+$signed( -{ 3'b0,x275 }<<<3'd2)+$signed( -{ 2'b0,x277 }<<<3'd1 )+$signed( { 1'b0,x278 }  )+$signed( -{ 2'b0,x279 }<<<3'd1 )+$signed( { 2'b0,x280 } <<<3'd1 )+$signed( { 2'b0,x282 } <<<3'd1 )+$signed( -{ 2'b0,x283 }<<<3'd1 )+$signed( { 1'b0,x284 }  )+$signed( -{ 2'b0,x286 }<<<3'd1 )+$signed( -{ 1'b0,x287 } )+$signed( -{ 3'b0,x288 }<<<3'd2)+$signed( -{ 2'b0,x289 }<<<3'd1 )+$signed( { 4'b0,x290 }<<<3'd3 )+$signed( { 3'b0,x292 }<<<3'd2 )+$signed( -{ 1'b0,x293 } )+$signed( -{ 2'b0,x294 }<<<3'd1 )+$signed( { 2'b0,x296 } <<<3'd1 )+$signed( { 1'b0,x297 }  )+$signed( -{ 2'b0,x298 }<<<3'd1 )+$signed( -{ 1'b0,x299 } )+$signed( { 2'b0,x300 } <<<3'd1 )+$signed( -{ 1'b0,x302 } )+$signed( { 2'b0,x303 } <<<3'd1 )+$signed( { 2'b0,x305 } <<<3'd1 )+$signed( { 3'b0,x306 }<<<3'd2 )+$signed( -{ 3'b0,x307 }<<<3'd2)+$signed( -{ 3'b0,x308 }<<<3'd2)+$signed( -{ 1'b0,x309 } )+$signed( -{ 3'b0,x311 }<<<3'd2)+$signed( -{ 2'b0,x312 }<<<3'd1 )+$signed( { 2'b0,x313 } <<<3'd1 )+$signed( -{ 3'b0,x314 }<<<3'd2)+$signed( { 2'b0,x315 } <<<3'd1 )+$signed( { 3'b0,x316 }<<<3'd2 )+$signed( { 3'b0,x317 }<<<3'd2 )+$signed( { 4'b0,x318 }<<<3'd3 )+$signed( { 3'b0,x319 }<<<3'd2 )+$signed( { 1'b0,x320 }  )+$signed( { 2'b0,x321 } <<<3'd1 )+$signed( -{ 1'b0,x323 } )+$signed( -{ 3'b0,x324 }<<<3'd2)+$signed( -{ 1'b0,x325 } )+$signed( -{ 2'b0,x327 }<<<3'd1 )+$signed( { 1'b0,x328 }  )+$signed( { 4'b0,x329 }<<<3'd3 )+$signed( { 1'b0,x330 }  )+$signed( { 3'b0,x331 }<<<3'd2 )+$signed( -{ 2'b0,x332 }<<<3'd1 )+$signed( -{ 2'b0,x333 }<<<3'd1 )+$signed( -{ 1'b0,x334 } )+$signed( { 2'b0,x335 } <<<3'd1 )+$signed( { 1'b0,x336 }  )+$signed( { 1'b0,x337 }  )+$signed( { 2'b0,x338 } <<<3'd1 )+$signed( -{ 3'b0,x339 }<<<3'd2)+$signed( { 1'b0,x340 }  )+$signed( { 3'b0,x342 }<<<3'd2 )+$signed( -{ 3'b0,x343 }<<<3'd2)+$signed( -{ 1'b0,x344 } )+$signed( -{ 3'b0,x345 }<<<3'd2)+$signed( { 2'b0,x346 } <<<3'd1 )+$signed( { 2'b0,x348 } <<<3'd1 )+$signed( -{ 3'b0,x349 }<<<3'd2)+$signed( { 2'b0,x351 } <<<3'd1 )+$signed( { 1'b0,x352 }  )+$signed( { 2'b0,x353 } <<<3'd1 )+$signed( { 2'b0,x354 } <<<3'd1 )+$signed( { 2'b0,x355 } <<<3'd1 )+$signed( { 2'b0,x357 } <<<3'd1 )+$signed( { 1'b0,x358 }  )+$signed( { 3'b0,x359 }<<<3'd2 )+$signed( { 2'b0,x360 } <<<3'd1 )+$signed( { 1'b0,x361 }  )+$signed( { 3'b0,x362 }<<<3'd2 )+$signed( { 2'b0,x363 } <<<3'd1 )+$signed( { 3'b0,x364 }<<<3'd2 )+$signed( { 1'b0,x365 }  )+$signed( -{ 3'b0,x366 }<<<3'd2)+$signed( -{ 2'b0,x368 }<<<3'd1 )+$signed( { 3'b0,x370 }<<<3'd2 )+$signed( { 3'b0,x372 }<<<3'd2 )+$signed( -{ 1'b0,x373 } )+$signed( { 3'b0,x374 }<<<3'd2 )+$signed( { 3'b0,x376 }<<<3'd2 )+$signed( { 1'b0,x377 }  )+$signed( { 2'b0,x378 } <<<3'd1 )+$signed( { 3'b0,x379 }<<<3'd2 )+$signed( { 1'b0,x380 }  )+$signed( { 4'b0,x381 }<<<3'd3 )+$signed( -{ 2'b0,x382 }<<<3'd1 )+$signed( { 1'b0,x383 }  )+$signed( -{ 2'b0,x384 }<<<3'd1 )+$signed( { 2'b0,x385 } <<<3'd1 )+$signed( -{ 2'b0,x386 }<<<3'd1 )+$signed( { 3'b0,x387 }<<<3'd2 )+$signed( -{ 2'b0,x388 }<<<3'd1 )+$signed( { 2'b0,x389 } <<<3'd1 )+$signed( { 3'b0,x390 }<<<3'd2 )+$signed( { 3'b0,x391 }<<<3'd2 )+$signed( -{ 2'b0,x392 }<<<3'd1 )+$signed( { 2'b0,x393 } <<<3'd1 )+$signed( -{ 1'b0,x394 } )+$signed( -{ 1'b0,x395 } )+$signed( -{ 2'b0,x396 }<<<3'd1 )+$signed( -{ 2'b0,x398 }<<<3'd1 )+$signed( { 3'b0,x400 }<<<3'd2 )+$signed( { 2'b0,x403 } <<<3'd1 )+$signed( -{ 3'b0,x404 }<<<3'd2)+$signed( { 1'b0,x405 }  )+$signed( -{ 2'b0,x406 }<<<3'd1 )+$signed( -{ 2'b0,x407 }<<<3'd1 )+$signed( { 3'b0,x408 }<<<3'd2 )+$signed( { 2'b0,x409 } <<<3'd1 )+$signed( { 3'b0,x410 }<<<3'd2 )+$signed( -{ 2'b0,x411 }<<<3'd1 )+$signed( { 2'b0,x412 } <<<3'd1 )+$signed( { 2'b0,x414 } <<<3'd1 )+$signed( -{ 1'b0,x416 } )+$signed( -{ 1'b0,x417 } )+$signed( { 2'b0,x418 } <<<3'd1 )+$signed( { 2'b0,x419 } <<<3'd1 )+$signed( -{ 1'b0,x420 } )+$signed( { 2'b0,x421 } <<<3'd1 )+$signed( -{ 2'b0,x422 }<<<3'd1 )+$signed( { 3'b0,x423 }<<<3'd2 )+$signed( { 3'b0,x425 }<<<3'd2 )+$signed( -{ 3'b0,x426 }<<<3'd2)+$signed( -{ 2'b0,x427 }<<<3'd1 )+$signed( -{ 3'b0,x428 }<<<3'd2)+$signed( -{ 2'b0,x429 }<<<3'd1 )+$signed( { 1'b0,x430 }  )+$signed( { 2'b0,x431 } <<<3'd1 )+$signed( { 1'b0,x432 }  )+$signed( { 2'b0,x433 } <<<3'd1 )+$signed( -{ 1'b0,x434 } )+$signed( -{ 2'b0,x436 }<<<3'd1 )+$signed( { 1'b0,x437 }  )+$signed( { 1'b0,x438 }  )+$signed( -{ 2'b0,x439 }<<<3'd1 )+$signed( -{ 2'b0,x442 }<<<3'd1 )+$signed( { 3'b0,x443 }<<<3'd2 )+$signed( { 1'b0,x444 }  )+$signed( { 2'b0,x445 } <<<3'd1 )+$signed( -{ 3'b0,x447 }<<<3'd2)+$signed( -{ 3'b0,x448 }<<<3'd2)+$signed( -{ 2'b0,x449 }<<<3'd1 )+$signed( { 2'b0,x451 } <<<3'd1 )+$signed( -{ 3'b0,x452 }<<<3'd2)+$signed( -{ 1'b0,x454 } )+$signed( -{ 2'b0,x455 }<<<3'd1 )+$signed( { 1'b0,x456 }  )+$signed( { 1'b0,x457 }  )+$signed( { 3'b0,x458 }<<<3'd2 )+$signed( { 3'b0,x459 }<<<3'd2 )+$signed( { 1'b0,x460 }  )+$signed( -{ 3'b0,x461 }<<<3'd2)+$signed( -{ 2'b0,x462 }<<<3'd1 )+$signed( -{ 2'b0,x463 }<<<3'd1 )+$signed( { 1'b0,x464 }  )+$signed( { 2'b0,x465 } <<<3'd1 )+$signed( -{ 3'b0,x466 }<<<3'd2)+$signed( { 1'b0,x467 }  )+$signed( { 2'b0,x468 } <<<3'd1 )+$signed( { 2'b0,x470 } <<<3'd1 )+$signed( { 3'b0,x471 }<<<3'd2 )+$signed( -{ 1'b0,x472 } )+$signed( -{ 2'b0,x473 }<<<3'd1 )+$signed( -{ 3'b0,x474 }<<<3'd2)+$signed( -{ 2'b0,x475 }<<<3'd1 )+$signed( { 1'b0,x476 }  )+$signed( -{ 3'b0,x480 }<<<3'd2)+$signed( { 2'b0,x481 } <<<3'd1 )+$signed( -{ 1'b0,x482 } )+$signed( -{ 3'b0,x483 }<<<3'd2)+$signed( { 3'b0,x484 }<<<3'd2 )+$signed( { 1'b0,x485 }  )+$signed( { 1'b0,x486 }  )+$signed( { 1'b0,x487 }  )+$signed( -{ 1'b0,x488 } )+$signed( { 1'b0,x489 }  )+$signed( { 1'b0,x490 }  )+$signed( -{ 3'b0,x491 }<<<3'd2)+$signed( -{ 1'b0,x492 } )+$signed( -{ 2'b0,x493 }<<<3'd1 )+$signed( { 2'b0,x495 } <<<3'd1 )-$signed(13'd24);
assign y3=temp_y[3][13] ==1'b1 ? 6'd0 :  
    temp_y[3][10] ==1'b1 ? 6'd63 : 
    temp_y[3][3]==1'b1 ? temp_y[3][9:4]+1'b1 : temp_y[3][9:4];
assign temp_y[4] = 
+$signed( { 2'b0,x0 } <<<3'd1 )+$signed( { 1'b0,x1 }  )+$signed( -{ 2'b0,x3 }<<<3'd1 )+$signed( -{ 1'b0,x4 } )+$signed( -{ 3'b0,x5 }<<<3'd2)+$signed( -{ 3'b0,x7 }<<<3'd2)+$signed( { 3'b0,x8 }<<<3'd2 )+$signed( -{ 4'b0, x9 }<<<3'd3 )+$signed( { 2'b0,x11 } <<<3'd1 )+$signed( -{ 3'b0,x12 }<<<3'd2)+$signed( { 3'b0,x13 }<<<3'd2 )+$signed( { 1'b0,x14 }  )+$signed( { 3'b0,x15 }<<<3'd2 )+$signed( { 3'b0,x16 }<<<3'd2 )+$signed( -{ 1'b0,x18 } )+$signed( { 3'b0,x19 }<<<3'd2 )+$signed( -{ 1'b0,x20 } )+$signed( -{ 1'b0,x22 } )+$signed( -{ 3'b0,x23 }<<<3'd2)+$signed( -{ 1'b0,x24 } )+$signed( -{ 3'b0,x25 }<<<3'd2)+$signed( { 2'b0,x26 } <<<3'd1 )+$signed( -{ 4'b0, x27 }<<<3'd3 )+$signed( { 1'b0,x28 }  )+$signed( { 1'b0,x29 }  )+$signed( { 1'b0,x30 }  )+$signed( { 2'b0,x31 } <<<3'd1 )+$signed( { 2'b0,x32 } <<<3'd1 )+$signed( { 1'b0,x33 }  )+$signed( { 1'b0,x34 }  )+$signed( -{ 1'b0,x35 } )+$signed( { 2'b0,x36 } <<<3'd1 )+$signed( { 3'b0,x37 }<<<3'd2 )+$signed( -{ 3'b0,x38 }<<<3'd2)+$signed( -{ 1'b0,x39 } )+$signed( -{ 2'b0,x40 }<<<3'd1 )+$signed( -{ 2'b0,x41 }<<<3'd1 )+$signed( { 1'b0,x43 }  )+$signed( { 2'b0,x44 } <<<3'd1 )+$signed( -{ 3'b0,x45 }<<<3'd2)+$signed( -{ 1'b0,x46 } )+$signed( { 1'b0,x47 }  )+$signed( { 1'b0,x48 }  )+$signed( { 2'b0,x49 } <<<3'd1 )+$signed( { 1'b0,x50 }  )+$signed( { 1'b0,x52 }  )+$signed( -{ 2'b0,x53 }<<<3'd1 )+$signed( { 3'b0,x55 }<<<3'd2 )+$signed( { 1'b0,x56 }  )+$signed( -{ 1'b0,x57 } )+$signed( { 2'b0,x58 } <<<3'd1 )+$signed( -{ 2'b0,x59 }<<<3'd1 )+$signed( { 3'b0,x61 }<<<3'd2 )+$signed( { 3'b0,x62 }<<<3'd2 )+$signed( -{ 3'b0,x63 }<<<3'd2)+$signed( { 3'b0,x64 }<<<3'd2 )+$signed( { 2'b0,x65 } <<<3'd1 )+$signed( { 2'b0,x67 } <<<3'd1 )+$signed( { 2'b0,x68 } <<<3'd1 )+$signed( { 2'b0,x69 } <<<3'd1 )+$signed( { 3'b0,x70 }<<<3'd2 )+$signed( { 3'b0,x71 }<<<3'd2 )+$signed( { 1'b0,x72 }  )+$signed( { 2'b0,x73 } <<<3'd1 )+$signed( -{ 1'b0,x74 } )+$signed( { 3'b0,x75 }<<<3'd2 )+$signed( { 1'b0,x76 }  )+$signed( -{ 2'b0,x77 }<<<3'd1 )+$signed( { 3'b0,x78 }<<<3'd2 )+$signed( -{ 2'b0,x79 }<<<3'd1 )+$signed( { 3'b0,x80 }<<<3'd2 )+$signed( -{ 3'b0,x81 }<<<3'd2)+$signed( { 2'b0,x84 } <<<3'd1 )+$signed( { 2'b0,x86 } <<<3'd1 )+$signed( -{ 1'b0,x87 } )+$signed( { 2'b0,x88 } <<<3'd1 )+$signed( -{ 1'b0,x89 } )+$signed( -{ 3'b0,x90 }<<<3'd2)+$signed( { 2'b0,x91 } <<<3'd1 )+$signed( -{ 2'b0,x92 }<<<3'd1 )+$signed( -{ 4'b0, x93 }<<<3'd3 )+$signed( { 3'b0,x95 }<<<3'd2 )+$signed( { 4'b0,x96 }<<<3'd3 )+$signed( { 3'b0,x97 }<<<3'd2 )+$signed( -{ 3'b0,x98 }<<<3'd2)+$signed( -{ 3'b0,x99 }<<<3'd2)+$signed( -{ 3'b0,x100 }<<<3'd2)+$signed( -{ 3'b0,x101 }<<<3'd2)+$signed( -{ 4'b0, x102 }<<<3'd3 )+$signed( { 1'b0,x103 }  )+$signed( { 3'b0,x104 }<<<3'd2 )+$signed( -{ 3'b0,x107 }<<<3'd2)+$signed( -{ 1'b0,x108 } )+$signed( -{ 2'b0,x109 }<<<3'd1 )+$signed( { 4'b0,x113 }<<<3'd3 )+$signed( { 3'b0,x114 }<<<3'd2 )+$signed( { 1'b0,x115 }  )+$signed( -{ 1'b0,x117 } )+$signed( { 1'b0,x118 }  )+$signed( -{ 2'b0,x119 }<<<3'd1 )+$signed( -{ 2'b0,x120 }<<<3'd1 )+$signed( { 2'b0,x121 } <<<3'd1 )+$signed( -{ 1'b0,x123 } )+$signed( -{ 2'b0,x124 }<<<3'd1 )+$signed( { 1'b0,x125 }  )+$signed( { 1'b0,x126 }  )+$signed( { 2'b0,x127 } <<<3'd1 )+$signed( -{ 1'b0,x128 } )+$signed( -{ 2'b0,x131 }<<<3'd1 )+$signed( { 1'b0,x132 }  )+$signed( { 3'b0,x133 }<<<3'd2 )+$signed( { 3'b0,x134 }<<<3'd2 )+$signed( -{ 3'b0,x135 }<<<3'd2)+$signed( -{ 2'b0,x136 }<<<3'd1 )+$signed( { 3'b0,x137 }<<<3'd2 )+$signed( { 2'b0,x139 } <<<3'd1 )+$signed( -{ 2'b0,x140 }<<<3'd1 )+$signed( { 2'b0,x141 } <<<3'd1 )+$signed( { 2'b0,x142 } <<<3'd1 )+$signed( -{ 2'b0,x143 }<<<3'd1 )+$signed( -{ 3'b0,x144 }<<<3'd2)+$signed( { 3'b0,x145 }<<<3'd2 )+$signed( { 1'b0,x146 }  )+$signed( { 2'b0,x147 } <<<3'd1 )+$signed( -{ 3'b0,x148 }<<<3'd2)+$signed( { 1'b0,x149 }  )+$signed( { 3'b0,x150 }<<<3'd2 )+$signed( -{ 3'b0,x151 }<<<3'd2)+$signed( { 2'b0,x152 } <<<3'd1 )+$signed( -{ 3'b0,x153 }<<<3'd2)+$signed( { 3'b0,x154 }<<<3'd2 )+$signed( { 3'b0,x156 }<<<3'd2 )+$signed( -{ 3'b0,x157 }<<<3'd2)+$signed( -{ 1'b0,x158 } )+$signed( -{ 3'b0,x159 }<<<3'd2)+$signed( -{ 2'b0,x160 }<<<3'd1 )+$signed( { 2'b0,x161 } <<<3'd1 )+$signed( -{ 1'b0,x162 } )+$signed( -{ 3'b0,x163 }<<<3'd2)+$signed( { 3'b0,x164 }<<<3'd2 )+$signed( -{ 2'b0,x166 }<<<3'd1 )+$signed( { 2'b0,x167 } <<<3'd1 )+$signed( { 3'b0,x168 }<<<3'd2 )+$signed( -{ 1'b0,x169 } )+$signed( { 2'b0,x170 } <<<3'd1 )+$signed( -{ 3'b0,x171 }<<<3'd2)+$signed( -{ 2'b0,x172 }<<<3'd1 )+$signed( -{ 3'b0,x175 }<<<3'd2)+$signed( -{ 3'b0,x176 }<<<3'd2)+$signed( { 1'b0,x177 }  )+$signed( -{ 3'b0,x178 }<<<3'd2)+$signed( -{ 3'b0,x179 }<<<3'd2)+$signed( { 3'b0,x180 }<<<3'd2 )+$signed( -{ 3'b0,x181 }<<<3'd2)+$signed( -{ 2'b0,x182 }<<<3'd1 )+$signed( -{ 2'b0,x183 }<<<3'd1 )+$signed( -{ 2'b0,x184 }<<<3'd1 )+$signed( { 2'b0,x185 } <<<3'd1 )+$signed( -{ 1'b0,x186 } )+$signed( -{ 3'b0,x187 }<<<3'd2)+$signed( { 2'b0,x188 } <<<3'd1 )+$signed( -{ 2'b0,x189 }<<<3'd1 )+$signed( { 2'b0,x190 } <<<3'd1 )+$signed( -{ 2'b0,x191 }<<<3'd1 )+$signed( -{ 2'b0,x192 }<<<3'd1 )+$signed( -{ 2'b0,x193 }<<<3'd1 )+$signed( -{ 1'b0,x194 } )+$signed( -{ 2'b0,x195 }<<<3'd1 )+$signed( { 1'b0,x196 }  )+$signed( -{ 3'b0,x197 }<<<3'd2)+$signed( -{ 2'b0,x198 }<<<3'd1 )+$signed( { 4'b0,x199 }<<<3'd3 )+$signed( { 3'b0,x200 }<<<3'd2 )+$signed( { 2'b0,x202 } <<<3'd1 )+$signed( { 3'b0,x203 }<<<3'd2 )+$signed( { 2'b0,x204 } <<<3'd1 )+$signed( { 3'b0,x205 }<<<3'd2 )+$signed( -{ 1'b0,x206 } )+$signed( -{ 3'b0,x207 }<<<3'd2)+$signed( { 1'b0,x208 }  )+$signed( -{ 1'b0,x209 } )+$signed( -{ 3'b0,x210 }<<<3'd2)+$signed( -{ 3'b0,x211 }<<<3'd2)+$signed( -{ 3'b0,x212 }<<<3'd2)+$signed( { 3'b0,x213 }<<<3'd2 )+$signed( -{ 3'b0,x214 }<<<3'd2)+$signed( -{ 2'b0,x215 }<<<3'd1 )+$signed( { 1'b0,x216 }  )+$signed( -{ 1'b0,x217 } )+$signed( { 1'b0,x218 }  )+$signed( { 2'b0,x219 } <<<3'd1 )+$signed( -{ 2'b0,x220 }<<<3'd1 )+$signed( { 1'b0,x221 }  )+$signed( { 3'b0,x222 }<<<3'd2 )+$signed( -{ 4'b0, x223 }<<<3'd3 )+$signed( { 2'b0,x224 } <<<3'd1 )+$signed( { 3'b0,x225 }<<<3'd2 )+$signed( -{ 1'b0,x226 } )+$signed( -{ 2'b0,x227 }<<<3'd1 )+$signed( -{ 2'b0,x228 }<<<3'd1 )+$signed( -{ 3'b0,x229 }<<<3'd2)+$signed( -{ 3'b0,x230 }<<<3'd2)+$signed( -{ 3'b0,x232 }<<<3'd2)+$signed( { 1'b0,x233 }  )+$signed( { 1'b0,x234 }  )+$signed( { 3'b0,x236 }<<<3'd2 )+$signed( -{ 2'b0,x237 }<<<3'd1 )+$signed( { 3'b0,x238 }<<<3'd2 )+$signed( -{ 2'b0,x239 }<<<3'd1 )+$signed( { 3'b0,x240 }<<<3'd2 )+$signed( -{ 2'b0,x241 }<<<3'd1 )+$signed( { 2'b0,x242 } <<<3'd1 )+$signed( -{ 1'b0,x243 } )+$signed( -{ 3'b0,x244 }<<<3'd2)+$signed( { 2'b0,x245 } <<<3'd1 )+$signed( -{ 2'b0,x246 }<<<3'd1 )+$signed( -{ 3'b0,x247 }<<<3'd2)+$signed( -{ 3'b0,x248 }<<<3'd2)+$signed( -{ 1'b0,x249 } )+$signed( -{ 1'b0,x250 } )+$signed( -{ 3'b0,x251 }<<<3'd2)+$signed( -{ 3'b0,x252 }<<<3'd2)+$signed( -{ 1'b0,x253 } )+$signed( { 1'b0,x254 }  )+$signed( -{ 2'b0,x256 }<<<3'd1 )+$signed( -{ 1'b0,x257 } )+$signed( { 3'b0,x258 }<<<3'd2 )+$signed( -{ 3'b0,x259 }<<<3'd2)+$signed( { 3'b0,x260 }<<<3'd2 )+$signed( -{ 3'b0,x261 }<<<3'd2)+$signed( { 3'b0,x262 }<<<3'd2 )+$signed( -{ 2'b0,x263 }<<<3'd1 )+$signed( -{ 2'b0,x264 }<<<3'd1 )+$signed( -{ 3'b0,x265 }<<<3'd2)+$signed( { 2'b0,x267 } <<<3'd1 )+$signed( -{ 4'b0, x268 }<<<3'd3 )+$signed( -{ 2'b0,x269 }<<<3'd1 )+$signed( -{ 3'b0,x271 }<<<3'd2)+$signed( { 3'b0,x272 }<<<3'd2 )+$signed( -{ 3'b0,x273 }<<<3'd2)+$signed( { 1'b0,x274 }  )+$signed( { 1'b0,x275 }  )+$signed( { 3'b0,x276 }<<<3'd2 )+$signed( -{ 1'b0,x277 } )+$signed( { 2'b0,x278 } <<<3'd1 )+$signed( -{ 2'b0,x279 }<<<3'd1 )+$signed( -{ 2'b0,x280 }<<<3'd1 )+$signed( -{ 2'b0,x281 }<<<3'd1 )+$signed( -{ 2'b0,x282 }<<<3'd1 )+$signed( -{ 4'b0, x283 }<<<3'd3 )+$signed( -{ 4'b0, x284 }<<<3'd3 )+$signed( { 2'b0,x285 } <<<3'd1 )+$signed( -{ 4'b0, x286 }<<<3'd3 )+$signed( -{ 2'b0,x287 }<<<3'd1 )+$signed( { 2'b0,x288 } <<<3'd1 )+$signed( -{ 1'b0,x290 } )+$signed( { 1'b0,x291 }  )+$signed( { 3'b0,x292 }<<<3'd2 )+$signed( { 1'b0,x293 }  )+$signed( { 2'b0,x294 } <<<3'd1 )+$signed( { 3'b0,x295 }<<<3'd2 )+$signed( { 2'b0,x296 } <<<3'd1 )+$signed( { 2'b0,x297 } <<<3'd1 )+$signed( -{ 1'b0,x298 } )+$signed( -{ 1'b0,x299 } )+$signed( -{ 1'b0,x300 } )+$signed( -{ 2'b0,x301 }<<<3'd1 )+$signed( { 2'b0,x302 } <<<3'd1 )+$signed( -{ 2'b0,x303 }<<<3'd1 )+$signed( { 3'b0,x304 }<<<3'd2 )+$signed( { 1'b0,x305 }  )+$signed( { 2'b0,x306 } <<<3'd1 )+$signed( { 2'b0,x307 } <<<3'd1 )+$signed( -{ 1'b0,x308 } )+$signed( { 3'b0,x310 }<<<3'd2 )+$signed( -{ 1'b0,x311 } )+$signed( -{ 2'b0,x312 }<<<3'd1 )+$signed( -{ 3'b0,x313 }<<<3'd2)+$signed( { 2'b0,x314 } <<<3'd1 )+$signed( { 2'b0,x315 } <<<3'd1 )+$signed( { 3'b0,x316 }<<<3'd2 )+$signed( { 1'b0,x317 }  )+$signed( -{ 4'b0, x318 }<<<3'd3 )+$signed( -{ 1'b0,x319 } )+$signed( { 2'b0,x320 } <<<3'd1 )+$signed( { 2'b0,x321 } <<<3'd1 )+$signed( -{ 2'b0,x322 }<<<3'd1 )+$signed( -{ 2'b0,x323 }<<<3'd1 )+$signed( { 2'b0,x324 } <<<3'd1 )+$signed( -{ 2'b0,x325 }<<<3'd1 )+$signed( { 2'b0,x327 } <<<3'd1 )+$signed( -{ 1'b0,x328 } )+$signed( { 3'b0,x330 }<<<3'd2 )+$signed( -{ 3'b0,x331 }<<<3'd2)+$signed( { 1'b0,x334 }  )+$signed( { 1'b0,x335 }  )+$signed( { 2'b0,x336 } <<<3'd1 )+$signed( { 1'b0,x338 }  )+$signed( -{ 3'b0,x339 }<<<3'd2)+$signed( -{ 1'b0,x340 } )+$signed( { 2'b0,x342 } <<<3'd1 )+$signed( { 4'b0,x343 }<<<3'd3 )+$signed( -{ 2'b0,x344 }<<<3'd1 )+$signed( { 3'b0,x345 }<<<3'd2 )+$signed( { 2'b0,x346 } <<<3'd1 )+$signed( { 2'b0,x347 } <<<3'd1 )+$signed( -{ 1'b0,x348 } )+$signed( { 2'b0,x349 } <<<3'd1 )+$signed( { 2'b0,x350 } <<<3'd1 )+$signed( -{ 2'b0,x351 }<<<3'd1 )+$signed( -{ 3'b0,x353 }<<<3'd2)+$signed( -{ 2'b0,x354 }<<<3'd1 )+$signed( -{ 2'b0,x355 }<<<3'd1 )+$signed( -{ 2'b0,x356 }<<<3'd1 )+$signed( -{ 2'b0,x357 }<<<3'd1 )+$signed( -{ 3'b0,x358 }<<<3'd2)+$signed( -{ 2'b0,x359 }<<<3'd1 )+$signed( { 3'b0,x361 }<<<3'd2 )+$signed( -{ 2'b0,x362 }<<<3'd1 )+$signed( { 3'b0,x364 }<<<3'd2 )+$signed( { 2'b0,x366 } <<<3'd1 )+$signed( { 3'b0,x368 }<<<3'd2 )+$signed( -{ 1'b0,x369 } )+$signed( -{ 3'b0,x370 }<<<3'd2)+$signed( { 2'b0,x371 } <<<3'd1 )+$signed( -{ 2'b0,x372 }<<<3'd1 )+$signed( -{ 1'b0,x373 } )+$signed( { 4'b0,x374 }<<<3'd3 )+$signed( -{ 1'b0,x375 } )+$signed( -{ 1'b0,x376 } )+$signed( -{ 2'b0,x377 }<<<3'd1 )+$signed( -{ 2'b0,x378 }<<<3'd1 )+$signed( { 1'b0,x379 }  )+$signed( { 2'b0,x380 } <<<3'd1 )+$signed( { 2'b0,x381 } <<<3'd1 )+$signed( { 3'b0,x382 }<<<3'd2 )+$signed( { 1'b0,x383 }  )+$signed( { 3'b0,x384 }<<<3'd2 )+$signed( -{ 2'b0,x386 }<<<3'd1 )+$signed( { 3'b0,x387 }<<<3'd2 )+$signed( { 1'b0,x388 }  )+$signed( -{ 2'b0,x389 }<<<3'd1 )+$signed( { 2'b0,x390 } <<<3'd1 )+$signed( -{ 4'b0, x391 }<<<3'd3 )+$signed( { 3'b0,x394 }<<<3'd2 )+$signed( -{ 3'b0,x395 }<<<3'd2)+$signed( -{ 2'b0,x396 }<<<3'd1 )+$signed( { 2'b0,x397 } <<<3'd1 )+$signed( -{ 2'b0,x399 }<<<3'd1 )+$signed( { 2'b0,x400 } <<<3'd1 )+$signed( { 2'b0,x401 } <<<3'd1 )+$signed( { 3'b0,x402 }<<<3'd2 )+$signed( -{ 2'b0,x403 }<<<3'd1 )+$signed( { 1'b0,x405 }  )+$signed( { 3'b0,x407 }<<<3'd2 )+$signed( -{ 1'b0,x408 } )+$signed( { 1'b0,x409 }  )+$signed( -{ 1'b0,x410 } )+$signed( -{ 1'b0,x411 } )+$signed( { 3'b0,x414 }<<<3'd2 )+$signed( { 3'b0,x415 }<<<3'd2 )+$signed( -{ 1'b0,x416 } )+$signed( { 3'b0,x418 }<<<3'd2 )+$signed( { 2'b0,x419 } <<<3'd1 )+$signed( { 3'b0,x420 }<<<3'd2 )+$signed( { 2'b0,x421 } <<<3'd1 )+$signed( { 1'b0,x422 }  )+$signed( { 2'b0,x423 } <<<3'd1 )+$signed( { 2'b0,x424 } <<<3'd1 )+$signed( -{ 1'b0,x425 } )+$signed( { 2'b0,x426 } <<<3'd1 )+$signed( { 1'b0,x427 }  )+$signed( -{ 2'b0,x428 }<<<3'd1 )+$signed( -{ 3'b0,x429 }<<<3'd2)+$signed( -{ 3'b0,x430 }<<<3'd2)+$signed( -{ 3'b0,x431 }<<<3'd2)+$signed( { 1'b0,x432 }  )+$signed( { 2'b0,x433 } <<<3'd1 )+$signed( { 2'b0,x435 } <<<3'd1 )+$signed( -{ 2'b0,x436 }<<<3'd1 )+$signed( { 2'b0,x437 } <<<3'd1 )+$signed( { 3'b0,x438 }<<<3'd2 )+$signed( { 3'b0,x439 }<<<3'd2 )+$signed( { 3'b0,x441 }<<<3'd2 )+$signed( { 1'b0,x442 }  )+$signed( -{ 2'b0,x443 }<<<3'd1 )+$signed( -{ 2'b0,x444 }<<<3'd1 )+$signed( -{ 2'b0,x446 }<<<3'd1 )+$signed( -{ 2'b0,x447 }<<<3'd1 )+$signed( -{ 3'b0,x449 }<<<3'd2)+$signed( -{ 1'b0,x450 } )+$signed( -{ 2'b0,x451 }<<<3'd1 )+$signed( -{ 2'b0,x452 }<<<3'd1 )+$signed( { 1'b0,x454 }  )+$signed( { 1'b0,x455 }  )+$signed( { 2'b0,x456 } <<<3'd1 )+$signed( -{ 3'b0,x457 }<<<3'd2)+$signed( -{ 3'b0,x458 }<<<3'd2)+$signed( -{ 1'b0,x460 } )+$signed( -{ 3'b0,x461 }<<<3'd2)+$signed( { 2'b0,x463 } <<<3'd1 )+$signed( -{ 2'b0,x464 }<<<3'd1 )+$signed( -{ 2'b0,x465 }<<<3'd1 )+$signed( -{ 1'b0,x466 } )+$signed( { 2'b0,x467 } <<<3'd1 )+$signed( -{ 4'b0, x468 }<<<3'd3 )+$signed( -{ 3'b0,x469 }<<<3'd2)+$signed( { 2'b0,x470 } <<<3'd1 )+$signed( -{ 1'b0,x472 } )+$signed( -{ 2'b0,x473 }<<<3'd1 )+$signed( -{ 3'b0,x474 }<<<3'd2)+$signed( { 2'b0,x475 } <<<3'd1 )+$signed( { 2'b0,x476 } <<<3'd1 )+$signed( -{ 3'b0,x478 }<<<3'd2)+$signed( { 3'b0,x479 }<<<3'd2 )+$signed( { 2'b0,x480 } <<<3'd1 )+$signed( { 3'b0,x481 }<<<3'd2 )+$signed( -{ 4'b0, x482 }<<<3'd3 )+$signed( -{ 2'b0,x483 }<<<3'd1 )+$signed( { 2'b0,x484 } <<<3'd1 )+$signed( -{ 2'b0,x487 }<<<3'd1 )+$signed( -{ 2'b0,x488 }<<<3'd1 )+$signed( { 1'b0,x489 }  )+$signed( { 1'b0,x490 }  )+$signed( -{ 3'b0,x491 }<<<3'd2)+$signed( { 2'b0,x492 } <<<3'd1 )+$signed( { 1'b0,x493 }  )+$signed( -{ 2'b0,x494 }<<<3'd1 )+$signed( -{ 1'b0,x495 } )+$signed(13'd8);
assign y4=temp_y[4][13] ==1'b1 ? 6'd0 :  
    temp_y[4][10] ==1'b1 ? 6'd63 : 
    temp_y[4][3]==1'b1 ? temp_y[4][9:4]+1'b1 : temp_y[4][9:4];
assign temp_y[5] = 
+$signed( { 2'b0,x0 } <<<3'd1 )+$signed( -{ 5'b0,x1 }<<<3'd4 )+$signed( -{ 3'b0,x2 }<<<3'd2)+$signed( -{ 3'b0,x3 }<<<3'd2)+$signed( { 3'b0,x4 }<<<3'd2 )+$signed( { 1'b0,x5 }  )+$signed( { 2'b0,x7 } <<<3'd1 )+$signed( { 1'b0,x8 }  )+$signed( -{ 3'b0,x10 }<<<3'd2)+$signed( -{ 3'b0,x11 }<<<3'd2)+$signed( { 1'b0,x12 }  )+$signed( -{ 2'b0,x13 }<<<3'd1 )+$signed( { 3'b0,x14 }<<<3'd2 )+$signed( { 1'b0,x15 }  )+$signed( -{ 2'b0,x16 }<<<3'd1 )+$signed( -{ 3'b0,x17 }<<<3'd2)+$signed( -{ 2'b0,x18 }<<<3'd1 )+$signed( { 3'b0,x19 }<<<3'd2 )+$signed( -{ 4'b0, x20 }<<<3'd3 )+$signed( { 3'b0,x21 }<<<3'd2 )+$signed( -{ 2'b0,x22 }<<<3'd1 )+$signed( { 2'b0,x24 } <<<3'd1 )+$signed( -{ 4'b0, x25 }<<<3'd3 )+$signed( { 1'b0,x26 }  )+$signed( { 3'b0,x27 }<<<3'd2 )+$signed( { 2'b0,x28 } <<<3'd1 )+$signed( { 3'b0,x29 }<<<3'd2 )+$signed( -{ 1'b0,x30 } )+$signed( -{ 1'b0,x31 } )+$signed( -{ 4'b0, x32 }<<<3'd3 )+$signed( { 1'b0,x33 }  )+$signed( { 1'b0,x35 }  )+$signed( { 3'b0,x36 }<<<3'd2 )+$signed( -{ 5'b0,x37 }<<<3'd4 )+$signed( -{ 2'b0,x39 }<<<3'd1 )+$signed( { 3'b0,x40 }<<<3'd2 )+$signed( -{ 3'b0,x41 }<<<3'd2)+$signed( { 3'b0,x42 }<<<3'd2 )+$signed( { 1'b0,x43 }  )+$signed( { 3'b0,x45 }<<<3'd2 )+$signed( -{ 5'b0,x47 }<<<3'd4 )+$signed( { 2'b0,x48 } <<<3'd1 )+$signed( { 3'b0,x49 }<<<3'd2 )+$signed( -{ 3'b0,x50 }<<<3'd2)+$signed( { 2'b0,x51 } <<<3'd1 )+$signed( -{ 2'b0,x52 }<<<3'd1 )+$signed( -{ 3'b0,x53 }<<<3'd2)+$signed( -{ 2'b0,x54 }<<<3'd1 )+$signed( -{ 5'b0,x55 }<<<3'd4 )+$signed( -{ 3'b0,x56 }<<<3'd2)+$signed( -{ 3'b0,x57 }<<<3'd2)+$signed( { 2'b0,x58 } <<<3'd1 )+$signed( -{ 2'b0,x59 }<<<3'd1 )+$signed( { 2'b0,x60 } <<<3'd1 )+$signed( -{ 3'b0,x63 }<<<3'd2)+$signed( -{ 3'b0,x64 }<<<3'd2)+$signed( -{ 5'b0,x65 }<<<3'd4 )+$signed( -{ 2'b0,x66 }<<<3'd1 )+$signed( -{ 3'b0,x67 }<<<3'd2)+$signed( -{ 4'b0, x68 }<<<3'd3 )+$signed( { 1'b0,x69 }  )+$signed( -{ 3'b0,x70 }<<<3'd2)+$signed( -{ 4'b0, x71 }<<<3'd3 )+$signed( { 2'b0,x72 } <<<3'd1 )+$signed( -{ 5'b0,x73 }<<<3'd4 )+$signed( { 1'b0,x74 }  )+$signed( { 1'b0,x77 }  )+$signed( -{ 1'b0,x79 } )+$signed( { 2'b0,x80 } <<<3'd1 )+$signed( { 1'b0,x82 }  )+$signed( { 2'b0,x83 } <<<3'd1 )+$signed( { 3'b0,x84 }<<<3'd2 )+$signed( -{ 2'b0,x85 }<<<3'd1 )+$signed( -{ 2'b0,x86 }<<<3'd1 )+$signed( { 2'b0,x87 } <<<3'd1 )+$signed( -{ 3'b0,x88 }<<<3'd2)+$signed( -{ 1'b0,x89 } )+$signed( { 2'b0,x90 } <<<3'd1 )+$signed( { 3'b0,x91 }<<<3'd2 )+$signed( -{ 3'b0,x92 }<<<3'd2)+$signed( { 3'b0,x93 }<<<3'd2 )+$signed( { 1'b0,x94 }  )+$signed( -{ 1'b0,x95 } )+$signed( { 1'b0,x96 }  )+$signed( -{ 3'b0,x97 }<<<3'd2)+$signed( { 4'b0,x98 }<<<3'd3 )+$signed( { 4'b0,x99 }<<<3'd3 )+$signed( { 1'b0,x100 }  )+$signed( -{ 4'b0, x102 }<<<3'd3 )+$signed( { 1'b0,x103 }  )+$signed( { 3'b0,x104 }<<<3'd2 )+$signed( { 1'b0,x108 }  )+$signed( { 3'b0,x109 }<<<3'd2 )+$signed( { 2'b0,x110 } <<<3'd1 )+$signed( { 2'b0,x111 } <<<3'd1 )+$signed( { 3'b0,x112 }<<<3'd2 )+$signed( { 2'b0,x113 } <<<3'd1 )+$signed( -{ 2'b0,x114 }<<<3'd1 )+$signed( { 3'b0,x115 }<<<3'd2 )+$signed( -{ 2'b0,x116 }<<<3'd1 )+$signed( -{ 3'b0,x117 }<<<3'd2)+$signed( { 3'b0,x118 }<<<3'd2 )+$signed( { 3'b0,x119 }<<<3'd2 )+$signed( -{ 3'b0,x121 }<<<3'd2)+$signed( -{ 4'b0, x122 }<<<3'd3 )+$signed( -{ 2'b0,x123 }<<<3'd1 )+$signed( { 1'b0,x124 }  )+$signed( -{ 2'b0,x125 }<<<3'd1 )+$signed( -{ 2'b0,x126 }<<<3'd1 )+$signed( -{ 5'b0,x127 }<<<3'd4 )+$signed( { 3'b0,x128 }<<<3'd2 )+$signed( -{ 3'b0,x129 }<<<3'd2)+$signed( { 2'b0,x130 } <<<3'd1 )+$signed( { 3'b0,x131 }<<<3'd2 )+$signed( -{ 1'b0,x132 } )+$signed( -{ 3'b0,x133 }<<<3'd2)+$signed( { 1'b0,x134 }  )+$signed( -{ 2'b0,x135 }<<<3'd1 )+$signed( { 3'b0,x137 }<<<3'd2 )+$signed( -{ 3'b0,x138 }<<<3'd2)+$signed( -{ 4'b0, x139 }<<<3'd3 )+$signed( -{ 1'b0,x140 } )+$signed( { 2'b0,x141 } <<<3'd1 )+$signed( -{ 3'b0,x143 }<<<3'd2)+$signed( -{ 3'b0,x144 }<<<3'd2)+$signed( -{ 3'b0,x145 }<<<3'd2)+$signed( -{ 1'b0,x146 } )+$signed( -{ 1'b0,x147 } )+$signed( { 3'b0,x148 }<<<3'd2 )+$signed( { 2'b0,x149 } <<<3'd1 )+$signed( { 2'b0,x150 } <<<3'd1 )+$signed( { 1'b0,x151 }  )+$signed( { 2'b0,x152 } <<<3'd1 )+$signed( -{ 1'b0,x153 } )+$signed( { 1'b0,x154 }  )+$signed( -{ 4'b0, x155 }<<<3'd3 )+$signed( { 3'b0,x156 }<<<3'd2 )+$signed( -{ 2'b0,x157 }<<<3'd1 )+$signed( -{ 1'b0,x158 } )+$signed( { 2'b0,x159 } <<<3'd1 )+$signed( -{ 4'b0, x160 }<<<3'd3 )+$signed( { 1'b0,x162 }  )+$signed( -{ 3'b0,x163 }<<<3'd2)+$signed( -{ 1'b0,x164 } )+$signed( -{ 4'b0, x165 }<<<3'd3 )+$signed( { 1'b0,x166 }  )+$signed( -{ 2'b0,x168 }<<<3'd1 )+$signed( { 2'b0,x169 } <<<3'd1 )+$signed( { 1'b0,x170 }  )+$signed( -{ 2'b0,x171 }<<<3'd1 )+$signed( -{ 2'b0,x172 }<<<3'd1 )+$signed( { 2'b0,x174 } <<<3'd1 )+$signed( -{ 3'b0,x177 }<<<3'd2)+$signed( { 2'b0,x178 } <<<3'd1 )+$signed( -{ 3'b0,x179 }<<<3'd2)+$signed( -{ 3'b0,x180 }<<<3'd2)+$signed( -{ 4'b0, x181 }<<<3'd3 )+$signed( -{ 1'b0,x182 } )+$signed( { 1'b0,x183 }  )+$signed( -{ 1'b0,x184 } )+$signed( -{ 1'b0,x185 } )+$signed( { 1'b0,x186 }  )+$signed( -{ 3'b0,x188 }<<<3'd2)+$signed( -{ 3'b0,x189 }<<<3'd2)+$signed( -{ 3'b0,x190 }<<<3'd2)+$signed( { 3'b0,x191 }<<<3'd2 )+$signed( { 1'b0,x192 }  )+$signed( { 2'b0,x193 } <<<3'd1 )+$signed( -{ 3'b0,x194 }<<<3'd2)+$signed( { 2'b0,x195 } <<<3'd1 )+$signed( -{ 1'b0,x196 } )+$signed( -{ 1'b0,x197 } )+$signed( -{ 3'b0,x198 }<<<3'd2)+$signed( -{ 5'b0,x199 }<<<3'd4 )+$signed( -{ 1'b0,x200 } )+$signed( { 3'b0,x201 }<<<3'd2 )+$signed( -{ 3'b0,x202 }<<<3'd2)+$signed( -{ 2'b0,x203 }<<<3'd1 )+$signed( -{ 1'b0,x205 } )+$signed( { 2'b0,x206 } <<<3'd1 )+$signed( -{ 3'b0,x207 }<<<3'd2)+$signed( { 1'b0,x210 }  )+$signed( { 1'b0,x211 }  )+$signed( { 2'b0,x212 } <<<3'd1 )+$signed( -{ 2'b0,x213 }<<<3'd1 )+$signed( -{ 1'b0,x214 } )+$signed( -{ 3'b0,x215 }<<<3'd2)+$signed( -{ 3'b0,x216 }<<<3'd2)+$signed( -{ 3'b0,x217 }<<<3'd2)+$signed( { 2'b0,x218 } <<<3'd1 )+$signed( -{ 3'b0,x219 }<<<3'd2)+$signed( { 3'b0,x220 }<<<3'd2 )+$signed( { 1'b0,x221 }  )+$signed( -{ 1'b0,x222 } )+$signed( { 2'b0,x223 } <<<3'd1 )+$signed( -{ 4'b0, x225 }<<<3'd3 )+$signed( -{ 3'b0,x226 }<<<3'd2)+$signed( -{ 2'b0,x227 }<<<3'd1 )+$signed( -{ 3'b0,x228 }<<<3'd2)+$signed( -{ 2'b0,x229 }<<<3'd1 )+$signed( { 4'b0,x230 }<<<3'd3 )+$signed( { 2'b0,x231 } <<<3'd1 )+$signed( { 3'b0,x232 }<<<3'd2 )+$signed( -{ 1'b0,x233 } )+$signed( -{ 2'b0,x234 }<<<3'd1 )+$signed( { 2'b0,x235 } <<<3'd1 )+$signed( -{ 2'b0,x236 }<<<3'd1 )+$signed( -{ 3'b0,x237 }<<<3'd2)+$signed( -{ 3'b0,x238 }<<<3'd2)+$signed( -{ 1'b0,x239 } )+$signed( -{ 3'b0,x240 }<<<3'd2)+$signed( { 2'b0,x241 } <<<3'd1 )+$signed( -{ 3'b0,x243 }<<<3'd2)+$signed( -{ 3'b0,x244 }<<<3'd2)+$signed( { 3'b0,x245 }<<<3'd2 )+$signed( { 3'b0,x246 }<<<3'd2 )+$signed( { 1'b0,x247 }  )+$signed( { 4'b0,x248 }<<<3'd3 )+$signed( -{ 2'b0,x249 }<<<3'd1 )+$signed( { 2'b0,x250 } <<<3'd1 )+$signed( { 3'b0,x251 }<<<3'd2 )+$signed( { 3'b0,x252 }<<<3'd2 )+$signed( -{ 4'b0, x253 }<<<3'd3 )+$signed( -{ 3'b0,x254 }<<<3'd2)+$signed( -{ 4'b0, x255 }<<<3'd3 )+$signed( -{ 3'b0,x256 }<<<3'd2)+$signed( -{ 2'b0,x257 }<<<3'd1 )+$signed( { 2'b0,x258 } <<<3'd1 )+$signed( { 3'b0,x259 }<<<3'd2 )+$signed( -{ 3'b0,x260 }<<<3'd2)+$signed( -{ 5'b0,x261 }<<<3'd4 )+$signed( -{ 3'b0,x262 }<<<3'd2)+$signed( { 2'b0,x263 } <<<3'd1 )+$signed( { 2'b0,x264 } <<<3'd1 )+$signed( { 2'b0,x265 } <<<3'd1 )+$signed( { 1'b0,x266 }  )+$signed( { 2'b0,x267 } <<<3'd1 )+$signed( { 2'b0,x268 } <<<3'd1 )+$signed( -{ 4'b0, x270 }<<<3'd3 )+$signed( -{ 3'b0,x271 }<<<3'd2)+$signed( { 3'b0,x272 }<<<3'd2 )+$signed( -{ 2'b0,x273 }<<<3'd1 )+$signed( -{ 2'b0,x274 }<<<3'd1 )+$signed( { 2'b0,x276 } <<<3'd1 )+$signed( { 4'b0,x277 }<<<3'd3 )+$signed( -{ 2'b0,x278 }<<<3'd1 )+$signed( -{ 2'b0,x279 }<<<3'd1 )+$signed( -{ 2'b0,x280 }<<<3'd1 )+$signed( { 3'b0,x281 }<<<3'd2 )+$signed( { 2'b0,x282 } <<<3'd1 )+$signed( -{ 1'b0,x283 } )+$signed( { 2'b0,x284 } <<<3'd1 )+$signed( -{ 3'b0,x286 }<<<3'd2)+$signed( { 1'b0,x287 }  )+$signed( { 3'b0,x288 }<<<3'd2 )+$signed( { 2'b0,x289 } <<<3'd1 )+$signed( { 2'b0,x290 } <<<3'd1 )+$signed( -{ 3'b0,x291 }<<<3'd2)+$signed( -{ 2'b0,x292 }<<<3'd1 )+$signed( -{ 4'b0, x293 }<<<3'd3 )+$signed( -{ 4'b0, x294 }<<<3'd3 )+$signed( -{ 4'b0, x296 }<<<3'd3 )+$signed( { 4'b0,x299 }<<<3'd3 )+$signed( -{ 3'b0,x300 }<<<3'd2)+$signed( -{ 2'b0,x301 }<<<3'd1 )+$signed( { 1'b0,x302 }  )+$signed( { 3'b0,x304 }<<<3'd2 )+$signed( { 1'b0,x305 }  )+$signed( { 3'b0,x307 }<<<3'd2 )+$signed( { 1'b0,x308 }  )+$signed( -{ 2'b0,x309 }<<<3'd1 )+$signed( { 2'b0,x310 } <<<3'd1 )+$signed( -{ 1'b0,x311 } )+$signed( -{ 3'b0,x312 }<<<3'd2)+$signed( { 3'b0,x313 }<<<3'd2 )+$signed( { 1'b0,x314 }  )+$signed( -{ 3'b0,x315 }<<<3'd2)+$signed( -{ 3'b0,x316 }<<<3'd2)+$signed( -{ 2'b0,x317 }<<<3'd1 )+$signed( -{ 4'b0, x318 }<<<3'd3 )+$signed( { 2'b0,x319 } <<<3'd1 )+$signed( -{ 4'b0, x321 }<<<3'd3 )+$signed( -{ 1'b0,x322 } )+$signed( -{ 2'b0,x323 }<<<3'd1 )+$signed( -{ 3'b0,x324 }<<<3'd2)+$signed( -{ 3'b0,x325 }<<<3'd2)+$signed( { 3'b0,x326 }<<<3'd2 )+$signed( -{ 2'b0,x327 }<<<3'd1 )+$signed( -{ 1'b0,x328 } )+$signed( { 1'b0,x329 }  )+$signed( -{ 2'b0,x330 }<<<3'd1 )+$signed( { 3'b0,x331 }<<<3'd2 )+$signed( -{ 2'b0,x333 }<<<3'd1 )+$signed( -{ 1'b0,x334 } )+$signed( { 2'b0,x335 } <<<3'd1 )+$signed( { 1'b0,x336 }  )+$signed( -{ 4'b0, x337 }<<<3'd3 )+$signed( { 3'b0,x338 }<<<3'd2 )+$signed( { 2'b0,x339 } <<<3'd1 )+$signed( { 1'b0,x341 }  )+$signed( -{ 2'b0,x343 }<<<3'd1 )+$signed( -{ 2'b0,x344 }<<<3'd1 )+$signed( { 2'b0,x345 } <<<3'd1 )+$signed( -{ 2'b0,x346 }<<<3'd1 )+$signed( { 3'b0,x347 }<<<3'd2 )+$signed( -{ 4'b0, x348 }<<<3'd3 )+$signed( { 2'b0,x349 } <<<3'd1 )+$signed( -{ 4'b0, x350 }<<<3'd3 )+$signed( { 3'b0,x351 }<<<3'd2 )+$signed( -{ 4'b0, x352 }<<<3'd3 )+$signed( { 1'b0,x353 }  )+$signed( -{ 1'b0,x354 } )+$signed( { 3'b0,x355 }<<<3'd2 )+$signed( -{ 1'b0,x356 } )+$signed( -{ 3'b0,x357 }<<<3'd2)+$signed( -{ 2'b0,x358 }<<<3'd1 )+$signed( -{ 1'b0,x359 } )+$signed( -{ 2'b0,x360 }<<<3'd1 )+$signed( -{ 1'b0,x361 } )+$signed( { 2'b0,x362 } <<<3'd1 )+$signed( { 3'b0,x363 }<<<3'd2 )+$signed( { 3'b0,x364 }<<<3'd2 )+$signed( { 3'b0,x365 }<<<3'd2 )+$signed( { 3'b0,x366 }<<<3'd2 )+$signed( { 3'b0,x368 }<<<3'd2 )+$signed( { 3'b0,x369 }<<<3'd2 )+$signed( { 4'b0,x370 }<<<3'd3 )+$signed( -{ 3'b0,x371 }<<<3'd2)+$signed( -{ 3'b0,x372 }<<<3'd2)+$signed( -{ 2'b0,x374 }<<<3'd1 )+$signed( -{ 2'b0,x375 }<<<3'd1 )+$signed( -{ 3'b0,x376 }<<<3'd2)+$signed( -{ 4'b0, x377 }<<<3'd3 )+$signed( { 5'b0,x378  }<<<3'd4 )+$signed( -{ 1'b0,x380 } )+$signed( -{ 3'b0,x381 }<<<3'd2)+$signed( { 3'b0,x382 }<<<3'd2 )+$signed( { 3'b0,x383 }<<<3'd2 )+$signed( { 3'b0,x384 }<<<3'd2 )+$signed( -{ 2'b0,x385 }<<<3'd1 )+$signed( { 1'b0,x386 }  )+$signed( { 3'b0,x387 }<<<3'd2 )+$signed( { 2'b0,x390 } <<<3'd1 )+$signed( { 3'b0,x392 }<<<3'd2 )+$signed( { 1'b0,x393 }  )+$signed( { 2'b0,x394 } <<<3'd1 )+$signed( -{ 2'b0,x396 }<<<3'd1 )+$signed( -{ 2'b0,x398 }<<<3'd1 )+$signed( { 2'b0,x400 } <<<3'd1 )+$signed( { 2'b0,x401 } <<<3'd1 )+$signed( -{ 2'b0,x402 }<<<3'd1 )+$signed( -{ 1'b0,x403 } )+$signed( { 2'b0,x404 } <<<3'd1 )+$signed( -{ 1'b0,x405 } )+$signed( -{ 2'b0,x406 }<<<3'd1 )+$signed( { 4'b0,x407 }<<<3'd3 )+$signed( -{ 2'b0,x408 }<<<3'd1 )+$signed( { 3'b0,x410 }<<<3'd2 )+$signed( -{ 3'b0,x411 }<<<3'd2)+$signed( { 1'b0,x412 }  )+$signed( { 1'b0,x414 }  )+$signed( { 3'b0,x415 }<<<3'd2 )+$signed( { 2'b0,x416 } <<<3'd1 )+$signed( { 3'b0,x417 }<<<3'd2 )+$signed( -{ 3'b0,x418 }<<<3'd2)+$signed( -{ 2'b0,x419 }<<<3'd1 )+$signed( { 4'b0,x420 }<<<3'd3 )+$signed( { 3'b0,x421 }<<<3'd2 )+$signed( -{ 1'b0,x422 } )+$signed( { 1'b0,x424 }  )+$signed( -{ 1'b0,x425 } )+$signed( { 3'b0,x426 }<<<3'd2 )+$signed( -{ 1'b0,x427 } )+$signed( -{ 2'b0,x428 }<<<3'd1 )+$signed( { 2'b0,x429 } <<<3'd1 )+$signed( -{ 2'b0,x430 }<<<3'd1 )+$signed( { 2'b0,x431 } <<<3'd1 )+$signed( -{ 3'b0,x432 }<<<3'd2)+$signed( { 4'b0,x433 }<<<3'd3 )+$signed( { 1'b0,x434 }  )+$signed( { 3'b0,x435 }<<<3'd2 )+$signed( -{ 3'b0,x436 }<<<3'd2)+$signed( -{ 3'b0,x438 }<<<3'd2)+$signed( { 1'b0,x439 }  )+$signed( -{ 1'b0,x440 } )+$signed( { 3'b0,x441 }<<<3'd2 )+$signed( { 2'b0,x442 } <<<3'd1 )+$signed( -{ 3'b0,x443 }<<<3'd2)+$signed( -{ 2'b0,x444 }<<<3'd1 )+$signed( { 3'b0,x445 }<<<3'd2 )+$signed( { 1'b0,x446 }  )+$signed( -{ 1'b0,x447 } )+$signed( -{ 2'b0,x448 }<<<3'd1 )+$signed( { 4'b0,x449 }<<<3'd3 )+$signed( -{ 2'b0,x450 }<<<3'd1 )+$signed( { 2'b0,x453 } <<<3'd1 )+$signed( -{ 3'b0,x454 }<<<3'd2)+$signed( { 2'b0,x455 } <<<3'd1 )+$signed( -{ 3'b0,x456 }<<<3'd2)+$signed( { 2'b0,x457 } <<<3'd1 )+$signed( { 3'b0,x458 }<<<3'd2 )+$signed( -{ 2'b0,x459 }<<<3'd1 )+$signed( { 4'b0,x460 }<<<3'd3 )+$signed( { 3'b0,x461 }<<<3'd2 )+$signed( { 3'b0,x462 }<<<3'd2 )+$signed( -{ 3'b0,x463 }<<<3'd2)+$signed( { 1'b0,x464 }  )+$signed( -{ 3'b0,x465 }<<<3'd2)+$signed( { 2'b0,x466 } <<<3'd1 )+$signed( -{ 4'b0, x467 }<<<3'd3 )+$signed( { 1'b0,x468 }  )+$signed( -{ 2'b0,x469 }<<<3'd1 )+$signed( { 3'b0,x470 }<<<3'd2 )+$signed( { 3'b0,x471 }<<<3'd2 )+$signed( -{ 4'b0, x472 }<<<3'd3 )+$signed( -{ 2'b0,x473 }<<<3'd1 )+$signed( { 2'b0,x475 } <<<3'd1 )+$signed( -{ 3'b0,x476 }<<<3'd2)+$signed( -{ 1'b0,x477 } )+$signed( { 4'b0,x478 }<<<3'd3 )+$signed( -{ 3'b0,x479 }<<<3'd2)+$signed( -{ 1'b0,x480 } )+$signed( -{ 5'b0,x481 }<<<3'd4 )+$signed( -{ 3'b0,x482 }<<<3'd2)+$signed( { 2'b0,x483 } <<<3'd1 )+$signed( -{ 2'b0,x484 }<<<3'd1 )+$signed( { 4'b0,x485 }<<<3'd3 )+$signed( { 4'b0,x487 }<<<3'd3 )+$signed( -{ 2'b0,x488 }<<<3'd1 )+$signed( { 1'b0,x489 }  )+$signed( { 1'b0,x490 }  )+$signed( { 2'b0,x491 } <<<3'd1 )+$signed( -{ 2'b0,x492 }<<<3'd1 )+$signed( -{ 2'b0,x493 }<<<3'd1 )+$signed( { 1'b0,x494 }  )+$signed( -{ 3'b0,x495 }<<<3'd2)-$signed(13'd16);
assign y5=temp_y[5][13] ==1'b1 ? 6'd0 :  
    temp_y[5][10] ==1'b1 ? 6'd63 : 
    temp_y[5][3]==1'b1 ? temp_y[5][9:4]+1'b1 : temp_y[5][9:4];
assign temp_y[6] = 
+$signed( -{ 3'b0,x0 }<<<3'd2)+$signed( { 3'b0,x1 }<<<3'd2 )+$signed( { 1'b0,x2 }  )+$signed( -{ 2'b0,x3 }<<<3'd1 )+$signed( -{ 2'b0,x5 }<<<3'd1 )+$signed( { 1'b0,x7 }  )+$signed( { 1'b0,x8 }  )+$signed( -{ 3'b0,x9 }<<<3'd2)+$signed( { 2'b0,x10 } <<<3'd1 )+$signed( { 3'b0,x11 }<<<3'd2 )+$signed( -{ 3'b0,x12 }<<<3'd2)+$signed( { 2'b0,x15 } <<<3'd1 )+$signed( { 1'b0,x17 }  )+$signed( -{ 1'b0,x18 } )+$signed( { 3'b0,x19 }<<<3'd2 )+$signed( { 2'b0,x20 } <<<3'd1 )+$signed( -{ 1'b0,x21 } )+$signed( -{ 2'b0,x23 }<<<3'd1 )+$signed( -{ 2'b0,x24 }<<<3'd1 )+$signed( -{ 3'b0,x25 }<<<3'd2)+$signed( { 1'b0,x26 }  )+$signed( -{ 2'b0,x27 }<<<3'd1 )+$signed( -{ 1'b0,x28 } )+$signed( { 2'b0,x29 } <<<3'd1 )+$signed( -{ 2'b0,x30 }<<<3'd1 )+$signed( { 3'b0,x31 }<<<3'd2 )+$signed( { 1'b0,x33 }  )+$signed( { 2'b0,x34 } <<<3'd1 )+$signed( -{ 2'b0,x36 }<<<3'd1 )+$signed( { 3'b0,x37 }<<<3'd2 )+$signed( { 3'b0,x38 }<<<3'd2 )+$signed( -{ 1'b0,x39 } )+$signed( { 3'b0,x40 }<<<3'd2 )+$signed( -{ 2'b0,x43 }<<<3'd1 )+$signed( { 3'b0,x44 }<<<3'd2 )+$signed( { 2'b0,x45 } <<<3'd1 )+$signed( { 2'b0,x46 } <<<3'd1 )+$signed( { 2'b0,x47 } <<<3'd1 )+$signed( { 1'b0,x48 }  )+$signed( { 3'b0,x49 }<<<3'd2 )+$signed( -{ 2'b0,x50 }<<<3'd1 )+$signed( { 2'b0,x51 } <<<3'd1 )+$signed( -{ 1'b0,x53 } )+$signed( { 1'b0,x54 }  )+$signed( { 3'b0,x55 }<<<3'd2 )+$signed( { 1'b0,x56 }  )+$signed( -{ 3'b0,x57 }<<<3'd2)+$signed( { 2'b0,x58 } <<<3'd1 )+$signed( -{ 2'b0,x59 }<<<3'd1 )+$signed( -{ 2'b0,x60 }<<<3'd1 )+$signed( -{ 1'b0,x61 } )+$signed( { 2'b0,x62 } <<<3'd1 )+$signed( -{ 3'b0,x63 }<<<3'd2)+$signed( { 2'b0,x64 } <<<3'd1 )+$signed( { 3'b0,x65 }<<<3'd2 )+$signed( { 1'b0,x66 }  )+$signed( -{ 1'b0,x67 } )+$signed( -{ 2'b0,x68 }<<<3'd1 )+$signed( { 2'b0,x69 } <<<3'd1 )+$signed( { 3'b0,x70 }<<<3'd2 )+$signed( { 2'b0,x71 } <<<3'd1 )+$signed( -{ 1'b0,x72 } )+$signed( { 1'b0,x73 }  )+$signed( { 1'b0,x74 }  )+$signed( -{ 4'b0, x75 }<<<3'd3 )+$signed( { 3'b0,x76 }<<<3'd2 )+$signed( -{ 2'b0,x77 }<<<3'd1 )+$signed( -{ 2'b0,x78 }<<<3'd1 )+$signed( { 2'b0,x79 } <<<3'd1 )+$signed( -{ 2'b0,x80 }<<<3'd1 )+$signed( -{ 3'b0,x81 }<<<3'd2)+$signed( -{ 1'b0,x82 } )+$signed( { 1'b0,x83 }  )+$signed( { 3'b0,x84 }<<<3'd2 )+$signed( { 2'b0,x86 } <<<3'd1 )+$signed( { 3'b0,x87 }<<<3'd2 )+$signed( -{ 1'b0,x89 } )+$signed( -{ 3'b0,x90 }<<<3'd2)+$signed( { 3'b0,x92 }<<<3'd2 )+$signed( { 1'b0,x93 }  )+$signed( { 3'b0,x94 }<<<3'd2 )+$signed( { 3'b0,x95 }<<<3'd2 )+$signed( { 3'b0,x96 }<<<3'd2 )+$signed( { 2'b0,x97 } <<<3'd1 )+$signed( { 1'b0,x98 }  )+$signed( { 2'b0,x99 } <<<3'd1 )+$signed( { 3'b0,x100 }<<<3'd2 )+$signed( -{ 1'b0,x101 } )+$signed( -{ 1'b0,x102 } )+$signed( { 1'b0,x103 }  )+$signed( { 1'b0,x104 }  )+$signed( { 3'b0,x105 }<<<3'd2 )+$signed( -{ 2'b0,x106 }<<<3'd1 )+$signed( { 1'b0,x107 }  )+$signed( -{ 3'b0,x108 }<<<3'd2)+$signed( -{ 2'b0,x109 }<<<3'd1 )+$signed( { 3'b0,x110 }<<<3'd2 )+$signed( { 4'b0,x111 }<<<3'd3 )+$signed( { 3'b0,x112 }<<<3'd2 )+$signed( { 1'b0,x113 }  )+$signed( { 1'b0,x114 }  )+$signed( -{ 1'b0,x115 } )+$signed( { 2'b0,x116 } <<<3'd1 )+$signed( { 1'b0,x117 }  )+$signed( { 3'b0,x118 }<<<3'd2 )+$signed( -{ 1'b0,x119 } )+$signed( -{ 1'b0,x120 } )+$signed( { 1'b0,x122 }  )+$signed( { 4'b0,x123 }<<<3'd3 )+$signed( -{ 3'b0,x124 }<<<3'd2)+$signed( { 2'b0,x125 } <<<3'd1 )+$signed( { 3'b0,x128 }<<<3'd2 )+$signed( -{ 3'b0,x129 }<<<3'd2)+$signed( -{ 1'b0,x130 } )+$signed( -{ 1'b0,x131 } )+$signed( -{ 2'b0,x132 }<<<3'd1 )+$signed( -{ 2'b0,x133 }<<<3'd1 )+$signed( { 1'b0,x134 }  )+$signed( -{ 1'b0,x135 } )+$signed( { 2'b0,x136 } <<<3'd1 )+$signed( -{ 2'b0,x137 }<<<3'd1 )+$signed( { 2'b0,x138 } <<<3'd1 )+$signed( { 2'b0,x139 } <<<3'd1 )+$signed( { 3'b0,x140 }<<<3'd2 )+$signed( { 2'b0,x141 } <<<3'd1 )+$signed( { 1'b0,x142 }  )+$signed( { 1'b0,x144 }  )+$signed( -{ 2'b0,x145 }<<<3'd1 )+$signed( { 2'b0,x146 } <<<3'd1 )+$signed( -{ 3'b0,x147 }<<<3'd2)+$signed( -{ 1'b0,x148 } )+$signed( -{ 1'b0,x149 } )+$signed( -{ 3'b0,x154 }<<<3'd2)+$signed( -{ 3'b0,x155 }<<<3'd2)+$signed( { 3'b0,x156 }<<<3'd2 )+$signed( { 2'b0,x157 } <<<3'd1 )+$signed( { 3'b0,x158 }<<<3'd2 )+$signed( { 3'b0,x159 }<<<3'd2 )+$signed( -{ 1'b0,x160 } )+$signed( { 1'b0,x161 }  )+$signed( { 1'b0,x162 }  )+$signed( -{ 1'b0,x163 } )+$signed( { 3'b0,x164 }<<<3'd2 )+$signed( { 3'b0,x165 }<<<3'd2 )+$signed( { 3'b0,x166 }<<<3'd2 )+$signed( { 1'b0,x167 }  )+$signed( -{ 2'b0,x168 }<<<3'd1 )+$signed( { 2'b0,x169 } <<<3'd1 )+$signed( { 3'b0,x170 }<<<3'd2 )+$signed( { 1'b0,x171 }  )+$signed( -{ 2'b0,x173 }<<<3'd1 )+$signed( { 3'b0,x174 }<<<3'd2 )+$signed( -{ 1'b0,x175 } )+$signed( -{ 1'b0,x176 } )+$signed( { 3'b0,x177 }<<<3'd2 )+$signed( -{ 2'b0,x178 }<<<3'd1 )+$signed( { 3'b0,x179 }<<<3'd2 )+$signed( { 3'b0,x180 }<<<3'd2 )+$signed( -{ 2'b0,x181 }<<<3'd1 )+$signed( { 3'b0,x182 }<<<3'd2 )+$signed( { 3'b0,x183 }<<<3'd2 )+$signed( { 2'b0,x184 } <<<3'd1 )+$signed( { 2'b0,x185 } <<<3'd1 )+$signed( -{ 3'b0,x186 }<<<3'd2)+$signed( -{ 1'b0,x189 } )+$signed( { 3'b0,x190 }<<<3'd2 )+$signed( -{ 3'b0,x191 }<<<3'd2)+$signed( { 3'b0,x192 }<<<3'd2 )+$signed( -{ 2'b0,x193 }<<<3'd1 )+$signed( { 1'b0,x194 }  )+$signed( { 3'b0,x195 }<<<3'd2 )+$signed( -{ 1'b0,x196 } )+$signed( { 3'b0,x197 }<<<3'd2 )+$signed( -{ 3'b0,x199 }<<<3'd2)+$signed( -{ 1'b0,x200 } )+$signed( -{ 2'b0,x201 }<<<3'd1 )+$signed( -{ 1'b0,x202 } )+$signed( { 2'b0,x205 } <<<3'd1 )+$signed( -{ 2'b0,x206 }<<<3'd1 )+$signed( { 2'b0,x207 } <<<3'd1 )+$signed( -{ 3'b0,x208 }<<<3'd2)+$signed( -{ 3'b0,x209 }<<<3'd2)+$signed( { 3'b0,x210 }<<<3'd2 )+$signed( { 1'b0,x211 }  )+$signed( { 3'b0,x212 }<<<3'd2 )+$signed( { 2'b0,x213 } <<<3'd1 )+$signed( { 1'b0,x215 }  )+$signed( -{ 4'b0, x217 }<<<3'd3 )+$signed( { 2'b0,x218 } <<<3'd1 )+$signed( -{ 3'b0,x220 }<<<3'd2)+$signed( -{ 1'b0,x221 } )+$signed( { 2'b0,x222 } <<<3'd1 )+$signed( { 2'b0,x223 } <<<3'd1 )+$signed( { 2'b0,x224 } <<<3'd1 )+$signed( -{ 2'b0,x225 }<<<3'd1 )+$signed( -{ 3'b0,x226 }<<<3'd2)+$signed( -{ 1'b0,x227 } )+$signed( { 1'b0,x229 }  )+$signed( -{ 2'b0,x231 }<<<3'd1 )+$signed( -{ 1'b0,x233 } )+$signed( { 1'b0,x234 }  )+$signed( -{ 2'b0,x235 }<<<3'd1 )+$signed( { 1'b0,x238 }  )+$signed( -{ 3'b0,x239 }<<<3'd2)+$signed( { 2'b0,x240 } <<<3'd1 )+$signed( { 4'b0,x241 }<<<3'd3 )+$signed( -{ 1'b0,x242 } )+$signed( -{ 2'b0,x243 }<<<3'd1 )+$signed( { 2'b0,x244 } <<<3'd1 )+$signed( { 3'b0,x245 }<<<3'd2 )+$signed( -{ 2'b0,x247 }<<<3'd1 )+$signed( { 1'b0,x248 }  )+$signed( -{ 1'b0,x250 } )+$signed( { 1'b0,x251 }  )+$signed( -{ 2'b0,x252 }<<<3'd1 )+$signed( -{ 2'b0,x253 }<<<3'd1 )+$signed( { 2'b0,x254 } <<<3'd1 )+$signed( { 3'b0,x255 }<<<3'd2 )+$signed( -{ 2'b0,x256 }<<<3'd1 )+$signed( -{ 2'b0,x257 }<<<3'd1 )+$signed( { 3'b0,x259 }<<<3'd2 )+$signed( { 1'b0,x260 }  )+$signed( -{ 3'b0,x261 }<<<3'd2)+$signed( { 2'b0,x262 } <<<3'd1 )+$signed( { 2'b0,x263 } <<<3'd1 )+$signed( -{ 2'b0,x264 }<<<3'd1 )+$signed( -{ 3'b0,x265 }<<<3'd2)+$signed( { 1'b0,x266 }  )+$signed( { 3'b0,x267 }<<<3'd2 )+$signed( { 2'b0,x268 } <<<3'd1 )+$signed( { 1'b0,x269 }  )+$signed( -{ 2'b0,x270 }<<<3'd1 )+$signed( -{ 3'b0,x271 }<<<3'd2)+$signed( -{ 2'b0,x272 }<<<3'd1 )+$signed( { 3'b0,x273 }<<<3'd2 )+$signed( -{ 3'b0,x274 }<<<3'd2)+$signed( -{ 2'b0,x275 }<<<3'd1 )+$signed( { 3'b0,x276 }<<<3'd2 )+$signed( { 3'b0,x277 }<<<3'd2 )+$signed( { 1'b0,x278 }  )+$signed( -{ 2'b0,x279 }<<<3'd1 )+$signed( -{ 4'b0, x280 }<<<3'd3 )+$signed( -{ 2'b0,x281 }<<<3'd1 )+$signed( { 3'b0,x282 }<<<3'd2 )+$signed( -{ 1'b0,x283 } )+$signed( { 1'b0,x284 }  )+$signed( { 2'b0,x285 } <<<3'd1 )+$signed( -{ 2'b0,x286 }<<<3'd1 )+$signed( -{ 2'b0,x287 }<<<3'd1 )+$signed( -{ 2'b0,x288 }<<<3'd1 )+$signed( { 1'b0,x289 }  )+$signed( -{ 2'b0,x290 }<<<3'd1 )+$signed( { 2'b0,x291 } <<<3'd1 )+$signed( -{ 1'b0,x292 } )+$signed( -{ 1'b0,x293 } )+$signed( { 1'b0,x294 }  )+$signed( -{ 3'b0,x295 }<<<3'd2)+$signed( -{ 1'b0,x296 } )+$signed( { 2'b0,x297 } <<<3'd1 )+$signed( { 2'b0,x298 } <<<3'd1 )+$signed( -{ 1'b0,x299 } )+$signed( { 1'b0,x300 }  )+$signed( { 1'b0,x302 }  )+$signed( -{ 3'b0,x303 }<<<3'd2)+$signed( { 3'b0,x304 }<<<3'd2 )+$signed( { 2'b0,x305 } <<<3'd1 )+$signed( { 1'b0,x307 }  )+$signed( -{ 3'b0,x308 }<<<3'd2)+$signed( -{ 2'b0,x309 }<<<3'd1 )+$signed( -{ 2'b0,x310 }<<<3'd1 )+$signed( { 4'b0,x311 }<<<3'd3 )+$signed( { 2'b0,x313 } <<<3'd1 )+$signed( { 1'b0,x314 }  )+$signed( -{ 2'b0,x315 }<<<3'd1 )+$signed( -{ 1'b0,x316 } )+$signed( { 2'b0,x317 } <<<3'd1 )+$signed( -{ 1'b0,x318 } )+$signed( { 3'b0,x320 }<<<3'd2 )+$signed( -{ 1'b0,x321 } )+$signed( { 2'b0,x322 } <<<3'd1 )+$signed( -{ 1'b0,x323 } )+$signed( { 3'b0,x324 }<<<3'd2 )+$signed( -{ 2'b0,x325 }<<<3'd1 )+$signed( { 3'b0,x326 }<<<3'd2 )+$signed( -{ 3'b0,x327 }<<<3'd2)+$signed( -{ 1'b0,x328 } )+$signed( -{ 2'b0,x329 }<<<3'd1 )+$signed( -{ 1'b0,x330 } )+$signed( -{ 2'b0,x331 }<<<3'd1 )+$signed( { 1'b0,x333 }  )+$signed( -{ 1'b0,x334 } )+$signed( { 3'b0,x336 }<<<3'd2 )+$signed( { 1'b0,x337 }  )+$signed( { 1'b0,x338 }  )+$signed( { 3'b0,x339 }<<<3'd2 )+$signed( { 2'b0,x340 } <<<3'd1 )+$signed( -{ 1'b0,x341 } )+$signed( { 1'b0,x342 }  )+$signed( -{ 3'b0,x344 }<<<3'd2)+$signed( { 2'b0,x345 } <<<3'd1 )+$signed( { 3'b0,x346 }<<<3'd2 )+$signed( -{ 3'b0,x347 }<<<3'd2)+$signed( -{ 2'b0,x348 }<<<3'd1 )+$signed( { 3'b0,x349 }<<<3'd2 )+$signed( { 3'b0,x350 }<<<3'd2 )+$signed( -{ 1'b0,x351 } )+$signed( { 2'b0,x352 } <<<3'd1 )+$signed( { 1'b0,x353 }  )+$signed( { 1'b0,x355 }  )+$signed( -{ 3'b0,x356 }<<<3'd2)+$signed( -{ 1'b0,x357 } )+$signed( -{ 1'b0,x358 } )+$signed( { 3'b0,x359 }<<<3'd2 )+$signed( -{ 3'b0,x360 }<<<3'd2)+$signed( { 2'b0,x361 } <<<3'd1 )+$signed( { 2'b0,x362 } <<<3'd1 )+$signed( { 3'b0,x363 }<<<3'd2 )+$signed( { 5'b0,x364  }<<<3'd4 )+$signed( { 3'b0,x365 }<<<3'd2 )+$signed( { 2'b0,x366 } <<<3'd1 )+$signed( -{ 1'b0,x367 } )+$signed( { 3'b0,x368 }<<<3'd2 )+$signed( -{ 3'b0,x369 }<<<3'd2)+$signed( { 1'b0,x370 }  )+$signed( { 2'b0,x372 } <<<3'd1 )+$signed( -{ 2'b0,x373 }<<<3'd1 )+$signed( { 3'b0,x374 }<<<3'd2 )+$signed( { 4'b0,x376 }<<<3'd3 )+$signed( { 3'b0,x377 }<<<3'd2 )+$signed( { 3'b0,x378 }<<<3'd2 )+$signed( -{ 2'b0,x379 }<<<3'd1 )+$signed( -{ 2'b0,x380 }<<<3'd1 )+$signed( { 3'b0,x381 }<<<3'd2 )+$signed( -{ 1'b0,x382 } )+$signed( -{ 3'b0,x383 }<<<3'd2)+$signed( { 2'b0,x384 } <<<3'd1 )+$signed( { 3'b0,x385 }<<<3'd2 )+$signed( -{ 3'b0,x386 }<<<3'd2)+$signed( { 3'b0,x387 }<<<3'd2 )+$signed( -{ 1'b0,x388 } )+$signed( { 3'b0,x389 }<<<3'd2 )+$signed( -{ 2'b0,x390 }<<<3'd1 )+$signed( { 2'b0,x391 } <<<3'd1 )+$signed( { 3'b0,x392 }<<<3'd2 )+$signed( -{ 2'b0,x393 }<<<3'd1 )+$signed( -{ 3'b0,x394 }<<<3'd2)+$signed( -{ 3'b0,x395 }<<<3'd2)+$signed( { 1'b0,x398 }  )+$signed( -{ 1'b0,x399 } )+$signed( { 3'b0,x400 }<<<3'd2 )+$signed( -{ 2'b0,x401 }<<<3'd1 )+$signed( -{ 2'b0,x403 }<<<3'd1 )+$signed( -{ 2'b0,x404 }<<<3'd1 )+$signed( { 2'b0,x405 } <<<3'd1 )+$signed( -{ 2'b0,x406 }<<<3'd1 )+$signed( { 2'b0,x407 } <<<3'd1 )+$signed( -{ 4'b0, x408 }<<<3'd3 )+$signed( -{ 2'b0,x409 }<<<3'd1 )+$signed( -{ 2'b0,x410 }<<<3'd1 )+$signed( { 3'b0,x411 }<<<3'd2 )+$signed( { 3'b0,x413 }<<<3'd2 )+$signed( { 1'b0,x414 }  )+$signed( { 3'b0,x415 }<<<3'd2 )+$signed( -{ 3'b0,x416 }<<<3'd2)+$signed( { 1'b0,x417 }  )+$signed( -{ 2'b0,x418 }<<<3'd1 )+$signed( { 3'b0,x420 }<<<3'd2 )+$signed( -{ 2'b0,x421 }<<<3'd1 )+$signed( -{ 3'b0,x422 }<<<3'd2)+$signed( { 2'b0,x423 } <<<3'd1 )+$signed( { 3'b0,x424 }<<<3'd2 )+$signed( { 3'b0,x426 }<<<3'd2 )+$signed( -{ 1'b0,x427 } )+$signed( { 3'b0,x428 }<<<3'd2 )+$signed( -{ 2'b0,x429 }<<<3'd1 )+$signed( { 2'b0,x430 } <<<3'd1 )+$signed( -{ 1'b0,x432 } )+$signed( { 1'b0,x433 }  )+$signed( -{ 3'b0,x435 }<<<3'd2)+$signed( -{ 1'b0,x436 } )+$signed( { 1'b0,x437 }  )+$signed( -{ 3'b0,x438 }<<<3'd2)+$signed( { 3'b0,x439 }<<<3'd2 )+$signed( { 1'b0,x440 }  )+$signed( { 3'b0,x441 }<<<3'd2 )+$signed( { 4'b0,x444 }<<<3'd3 )+$signed( -{ 1'b0,x445 } )+$signed( -{ 4'b0, x446 }<<<3'd3 )+$signed( { 2'b0,x447 } <<<3'd1 )+$signed( { 1'b0,x448 }  )+$signed( { 1'b0,x449 }  )+$signed( { 2'b0,x450 } <<<3'd1 )+$signed( { 3'b0,x452 }<<<3'd2 )+$signed( -{ 2'b0,x453 }<<<3'd1 )+$signed( -{ 1'b0,x454 } )+$signed( { 2'b0,x455 } <<<3'd1 )+$signed( -{ 3'b0,x456 }<<<3'd2)+$signed( { 3'b0,x457 }<<<3'd2 )+$signed( { 3'b0,x459 }<<<3'd2 )+$signed( -{ 1'b0,x460 } )+$signed( -{ 3'b0,x461 }<<<3'd2)+$signed( -{ 1'b0,x462 } )+$signed( -{ 1'b0,x463 } )+$signed( { 3'b0,x464 }<<<3'd2 )+$signed( { 2'b0,x465 } <<<3'd1 )+$signed( -{ 2'b0,x466 }<<<3'd1 )+$signed( { 2'b0,x467 } <<<3'd1 )+$signed( { 4'b0,x468 }<<<3'd3 )+$signed( -{ 2'b0,x470 }<<<3'd1 )+$signed( { 2'b0,x471 } <<<3'd1 )+$signed( -{ 1'b0,x472 } )+$signed( { 3'b0,x473 }<<<3'd2 )+$signed( { 1'b0,x474 }  )+$signed( { 1'b0,x475 }  )+$signed( { 2'b0,x476 } <<<3'd1 )+$signed( { 3'b0,x477 }<<<3'd2 )+$signed( { 3'b0,x478 }<<<3'd2 )+$signed( -{ 1'b0,x479 } )+$signed( { 1'b0,x480 }  )+$signed( { 3'b0,x481 }<<<3'd2 )+$signed( { 1'b0,x482 }  )+$signed( { 3'b0,x483 }<<<3'd2 )+$signed( { 1'b0,x484 }  )+$signed( -{ 3'b0,x485 }<<<3'd2)+$signed( { 2'b0,x486 } <<<3'd1 )+$signed( -{ 2'b0,x487 }<<<3'd1 )+$signed( { 1'b0,x488 }  )+$signed( { 3'b0,x490 }<<<3'd2 )+$signed( { 1'b0,x492 }  )+$signed( { 2'b0,x493 } <<<3'd1 )+$signed( { 3'b0,x494 }<<<3'd2 )+$signed( -{ 2'b0,x495 }<<<3'd1 )-$signed(13'd48);
assign y6=temp_y[6][13] ==1'b1 ? 6'd0 :  
    temp_y[6][10] ==1'b1 ? 6'd63 : 
    temp_y[6][3]==1'b1 ? temp_y[6][9:4]+1'b1 : temp_y[6][9:4];
assign temp_y[7] = 
+$signed( -{ 1'b0,x0 } )+$signed( -{ 2'b0,x1 }<<<3'd1 )+$signed( -{ 2'b0,x3 }<<<3'd1 )+$signed( -{ 3'b0,x5 }<<<3'd2)+$signed( { 3'b0,x6 }<<<3'd2 )+$signed( { 4'b0,x7 }<<<3'd3 )+$signed( { 3'b0,x8 }<<<3'd2 )+$signed( -{ 1'b0,x9 } )+$signed( -{ 1'b0,x10 } )+$signed( -{ 3'b0,x12 }<<<3'd2)+$signed( -{ 2'b0,x13 }<<<3'd1 )+$signed( -{ 2'b0,x14 }<<<3'd1 )+$signed( { 3'b0,x15 }<<<3'd2 )+$signed( -{ 1'b0,x17 } )+$signed( -{ 2'b0,x19 }<<<3'd1 )+$signed( -{ 3'b0,x20 }<<<3'd2)+$signed( -{ 3'b0,x21 }<<<3'd2)+$signed( { 2'b0,x22 } <<<3'd1 )+$signed( -{ 1'b0,x23 } )+$signed( -{ 1'b0,x24 } )+$signed( { 3'b0,x25 }<<<3'd2 )+$signed( { 3'b0,x26 }<<<3'd2 )+$signed( -{ 1'b0,x27 } )+$signed( -{ 1'b0,x28 } )+$signed( { 2'b0,x29 } <<<3'd1 )+$signed( { 1'b0,x30 }  )+$signed( { 1'b0,x31 }  )+$signed( { 2'b0,x33 } <<<3'd1 )+$signed( { 1'b0,x34 }  )+$signed( -{ 1'b0,x35 } )+$signed( -{ 2'b0,x36 }<<<3'd1 )+$signed( -{ 2'b0,x37 }<<<3'd1 )+$signed( -{ 1'b0,x38 } )+$signed( -{ 2'b0,x39 }<<<3'd1 )+$signed( { 2'b0,x40 } <<<3'd1 )+$signed( { 2'b0,x41 } <<<3'd1 )+$signed( { 2'b0,x42 } <<<3'd1 )+$signed( { 3'b0,x43 }<<<3'd2 )+$signed( { 2'b0,x44 } <<<3'd1 )+$signed( -{ 1'b0,x45 } )+$signed( { 2'b0,x46 } <<<3'd1 )+$signed( { 2'b0,x48 } <<<3'd1 )+$signed( { 2'b0,x49 } <<<3'd1 )+$signed( { 3'b0,x50 }<<<3'd2 )+$signed( -{ 2'b0,x52 }<<<3'd1 )+$signed( { 1'b0,x54 }  )+$signed( -{ 2'b0,x56 }<<<3'd1 )+$signed( -{ 1'b0,x57 } )+$signed( { 2'b0,x58 } <<<3'd1 )+$signed( -{ 2'b0,x59 }<<<3'd1 )+$signed( { 1'b0,x60 }  )+$signed( { 3'b0,x61 }<<<3'd2 )+$signed( { 3'b0,x62 }<<<3'd2 )+$signed( -{ 2'b0,x63 }<<<3'd1 )+$signed( { 1'b0,x65 }  )+$signed( -{ 2'b0,x66 }<<<3'd1 )+$signed( -{ 2'b0,x67 }<<<3'd1 )+$signed( { 1'b0,x68 }  )+$signed( { 3'b0,x69 }<<<3'd2 )+$signed( { 1'b0,x70 }  )+$signed( -{ 2'b0,x71 }<<<3'd1 )+$signed( { 1'b0,x72 }  )+$signed( -{ 3'b0,x75 }<<<3'd2)+$signed( { 3'b0,x76 }<<<3'd2 )+$signed( { 1'b0,x77 }  )+$signed( -{ 1'b0,x78 } )+$signed( { 3'b0,x79 }<<<3'd2 )+$signed( { 2'b0,x80 } <<<3'd1 )+$signed( { 3'b0,x81 }<<<3'd2 )+$signed( { 2'b0,x83 } <<<3'd1 )+$signed( -{ 2'b0,x84 }<<<3'd1 )+$signed( -{ 2'b0,x86 }<<<3'd1 )+$signed( { 2'b0,x87 } <<<3'd1 )+$signed( -{ 2'b0,x89 }<<<3'd1 )+$signed( { 2'b0,x90 } <<<3'd1 )+$signed( -{ 2'b0,x91 }<<<3'd1 )+$signed( -{ 3'b0,x93 }<<<3'd2)+$signed( -{ 1'b0,x94 } )+$signed( -{ 1'b0,x95 } )+$signed( { 3'b0,x96 }<<<3'd2 )+$signed( { 3'b0,x98 }<<<3'd2 )+$signed( -{ 2'b0,x99 }<<<3'd1 )+$signed( { 3'b0,x100 }<<<3'd2 )+$signed( -{ 1'b0,x101 } )+$signed( { 2'b0,x103 } <<<3'd1 )+$signed( { 2'b0,x104 } <<<3'd1 )+$signed( { 1'b0,x105 }  )+$signed( { 1'b0,x106 }  )+$signed( -{ 2'b0,x107 }<<<3'd1 )+$signed( -{ 2'b0,x108 }<<<3'd1 )+$signed( -{ 2'b0,x109 }<<<3'd1 )+$signed( { 2'b0,x110 } <<<3'd1 )+$signed( { 3'b0,x111 }<<<3'd2 )+$signed( -{ 3'b0,x112 }<<<3'd2)+$signed( { 1'b0,x113 }  )+$signed( { 2'b0,x114 } <<<3'd1 )+$signed( { 3'b0,x116 }<<<3'd2 )+$signed( -{ 3'b0,x117 }<<<3'd2)+$signed( { 3'b0,x118 }<<<3'd2 )+$signed( -{ 2'b0,x119 }<<<3'd1 )+$signed( { 2'b0,x121 } <<<3'd1 )+$signed( { 3'b0,x122 }<<<3'd2 )+$signed( { 1'b0,x125 }  )+$signed( -{ 2'b0,x127 }<<<3'd1 )+$signed( { 2'b0,x128 } <<<3'd1 )+$signed( -{ 1'b0,x129 } )+$signed( { 1'b0,x130 }  )+$signed( -{ 1'b0,x131 } )+$signed( -{ 1'b0,x132 } )+$signed( { 1'b0,x133 }  )+$signed( { 2'b0,x134 } <<<3'd1 )+$signed( { 3'b0,x135 }<<<3'd2 )+$signed( { 3'b0,x136 }<<<3'd2 )+$signed( -{ 3'b0,x137 }<<<3'd2)+$signed( -{ 2'b0,x138 }<<<3'd1 )+$signed( { 2'b0,x139 } <<<3'd1 )+$signed( -{ 2'b0,x140 }<<<3'd1 )+$signed( { 3'b0,x141 }<<<3'd2 )+$signed( -{ 2'b0,x143 }<<<3'd1 )+$signed( -{ 2'b0,x144 }<<<3'd1 )+$signed( { 1'b0,x145 }  )+$signed( -{ 2'b0,x147 }<<<3'd1 )+$signed( { 2'b0,x148 } <<<3'd1 )+$signed( { 2'b0,x149 } <<<3'd1 )+$signed( -{ 2'b0,x150 }<<<3'd1 )+$signed( { 2'b0,x152 } <<<3'd1 )+$signed( { 3'b0,x153 }<<<3'd2 )+$signed( { 2'b0,x154 } <<<3'd1 )+$signed( { 3'b0,x156 }<<<3'd2 )+$signed( -{ 2'b0,x157 }<<<3'd1 )+$signed( { 1'b0,x158 }  )+$signed( { 3'b0,x159 }<<<3'd2 )+$signed( -{ 2'b0,x161 }<<<3'd1 )+$signed( -{ 3'b0,x162 }<<<3'd2)+$signed( { 2'b0,x163 } <<<3'd1 )+$signed( { 2'b0,x164 } <<<3'd1 )+$signed( -{ 1'b0,x165 } )+$signed( { 3'b0,x166 }<<<3'd2 )+$signed( { 3'b0,x167 }<<<3'd2 )+$signed( { 3'b0,x168 }<<<3'd2 )+$signed( { 3'b0,x169 }<<<3'd2 )+$signed( -{ 3'b0,x170 }<<<3'd2)+$signed( { 1'b0,x171 }  )+$signed( { 2'b0,x172 } <<<3'd1 )+$signed( { 2'b0,x173 } <<<3'd1 )+$signed( -{ 2'b0,x175 }<<<3'd1 )+$signed( -{ 2'b0,x176 }<<<3'd1 )+$signed( { 1'b0,x177 }  )+$signed( -{ 1'b0,x178 } )+$signed( { 3'b0,x179 }<<<3'd2 )+$signed( -{ 2'b0,x180 }<<<3'd1 )+$signed( { 1'b0,x183 }  )+$signed( { 3'b0,x184 }<<<3'd2 )+$signed( { 2'b0,x185 } <<<3'd1 )+$signed( { 3'b0,x186 }<<<3'd2 )+$signed( -{ 3'b0,x188 }<<<3'd2)+$signed( -{ 1'b0,x189 } )+$signed( { 3'b0,x191 }<<<3'd2 )+$signed( -{ 2'b0,x193 }<<<3'd1 )+$signed( -{ 3'b0,x194 }<<<3'd2)+$signed( { 3'b0,x196 }<<<3'd2 )+$signed( { 3'b0,x197 }<<<3'd2 )+$signed( -{ 1'b0,x198 } )+$signed( -{ 1'b0,x199 } )+$signed( { 2'b0,x200 } <<<3'd1 )+$signed( -{ 4'b0, x201 }<<<3'd3 )+$signed( { 2'b0,x202 } <<<3'd1 )+$signed( { 1'b0,x203 }  )+$signed( -{ 1'b0,x204 } )+$signed( { 3'b0,x205 }<<<3'd2 )+$signed( { 2'b0,x206 } <<<3'd1 )+$signed( { 3'b0,x207 }<<<3'd2 )+$signed( { 2'b0,x209 } <<<3'd1 )+$signed( -{ 2'b0,x210 }<<<3'd1 )+$signed( { 2'b0,x211 } <<<3'd1 )+$signed( -{ 2'b0,x212 }<<<3'd1 )+$signed( { 3'b0,x214 }<<<3'd2 )+$signed( -{ 2'b0,x215 }<<<3'd1 )+$signed( -{ 1'b0,x216 } )+$signed( -{ 1'b0,x217 } )+$signed( { 1'b0,x218 }  )+$signed( { 2'b0,x219 } <<<3'd1 )+$signed( -{ 2'b0,x220 }<<<3'd1 )+$signed( -{ 1'b0,x221 } )+$signed( { 1'b0,x222 }  )+$signed( -{ 2'b0,x223 }<<<3'd1 )+$signed( { 3'b0,x224 }<<<3'd2 )+$signed( { 2'b0,x225 } <<<3'd1 )+$signed( { 3'b0,x226 }<<<3'd2 )+$signed( { 2'b0,x227 } <<<3'd1 )+$signed( -{ 3'b0,x228 }<<<3'd2)+$signed( -{ 3'b0,x229 }<<<3'd2)+$signed( -{ 3'b0,x230 }<<<3'd2)+$signed( -{ 1'b0,x233 } )+$signed( { 2'b0,x234 } <<<3'd1 )+$signed( -{ 1'b0,x235 } )+$signed( { 1'b0,x237 }  )+$signed( { 2'b0,x238 } <<<3'd1 )+$signed( -{ 1'b0,x240 } )+$signed( { 2'b0,x241 } <<<3'd1 )+$signed( -{ 2'b0,x242 }<<<3'd1 )+$signed( { 1'b0,x243 }  )+$signed( { 2'b0,x244 } <<<3'd1 )+$signed( { 3'b0,x245 }<<<3'd2 )+$signed( { 1'b0,x246 }  )+$signed( { 3'b0,x247 }<<<3'd2 )+$signed( { 3'b0,x248 }<<<3'd2 )+$signed( { 4'b0,x250 }<<<3'd3 )+$signed( { 2'b0,x252 } <<<3'd1 )+$signed( -{ 2'b0,x253 }<<<3'd1 )+$signed( -{ 1'b0,x254 } )+$signed( { 2'b0,x255 } <<<3'd1 )+$signed( -{ 3'b0,x256 }<<<3'd2)+$signed( -{ 1'b0,x257 } )+$signed( { 3'b0,x259 }<<<3'd2 )+$signed( -{ 1'b0,x260 } )+$signed( -{ 3'b0,x261 }<<<3'd2)+$signed( -{ 1'b0,x262 } )+$signed( { 3'b0,x263 }<<<3'd2 )+$signed( -{ 1'b0,x264 } )+$signed( { 2'b0,x265 } <<<3'd1 )+$signed( { 3'b0,x266 }<<<3'd2 )+$signed( { 3'b0,x267 }<<<3'd2 )+$signed( -{ 1'b0,x268 } )+$signed( { 1'b0,x269 }  )+$signed( { 3'b0,x270 }<<<3'd2 )+$signed( -{ 2'b0,x271 }<<<3'd1 )+$signed( -{ 2'b0,x272 }<<<3'd1 )+$signed( { 2'b0,x274 } <<<3'd1 )+$signed( { 1'b0,x275 }  )+$signed( { 2'b0,x276 } <<<3'd1 )+$signed( { 2'b0,x277 } <<<3'd1 )+$signed( { 3'b0,x278 }<<<3'd2 )+$signed( { 1'b0,x279 }  )+$signed( { 3'b0,x280 }<<<3'd2 )+$signed( { 3'b0,x281 }<<<3'd2 )+$signed( -{ 2'b0,x282 }<<<3'd1 )+$signed( -{ 1'b0,x283 } )+$signed( -{ 2'b0,x285 }<<<3'd1 )+$signed( -{ 4'b0, x286 }<<<3'd3 )+$signed( { 1'b0,x287 }  )+$signed( { 1'b0,x288 }  )+$signed( { 2'b0,x289 } <<<3'd1 )+$signed( -{ 1'b0,x290 } )+$signed( -{ 1'b0,x291 } )+$signed( -{ 3'b0,x292 }<<<3'd2)+$signed( -{ 3'b0,x293 }<<<3'd2)+$signed( { 3'b0,x294 }<<<3'd2 )+$signed( { 3'b0,x295 }<<<3'd2 )+$signed( { 3'b0,x296 }<<<3'd2 )+$signed( { 1'b0,x297 }  )+$signed( { 1'b0,x298 }  )+$signed( { 1'b0,x299 }  )+$signed( { 2'b0,x300 } <<<3'd1 )+$signed( { 1'b0,x301 }  )+$signed( -{ 2'b0,x302 }<<<3'd1 )+$signed( -{ 4'b0, x303 }<<<3'd3 )+$signed( -{ 2'b0,x304 }<<<3'd1 )+$signed( -{ 4'b0, x305 }<<<3'd3 )+$signed( { 2'b0,x306 } <<<3'd1 )+$signed( -{ 1'b0,x308 } )+$signed( -{ 1'b0,x310 } )+$signed( { 1'b0,x311 }  )+$signed( -{ 2'b0,x312 }<<<3'd1 )+$signed( { 2'b0,x313 } <<<3'd1 )+$signed( -{ 1'b0,x315 } )+$signed( -{ 1'b0,x316 } )+$signed( { 4'b0,x317 }<<<3'd3 )+$signed( { 2'b0,x319 } <<<3'd1 )+$signed( { 3'b0,x320 }<<<3'd2 )+$signed( { 3'b0,x321 }<<<3'd2 )+$signed( -{ 2'b0,x322 }<<<3'd1 )+$signed( -{ 2'b0,x323 }<<<3'd1 )+$signed( { 1'b0,x324 }  )+$signed( -{ 1'b0,x325 } )+$signed( -{ 3'b0,x327 }<<<3'd2)+$signed( -{ 1'b0,x328 } )+$signed( -{ 2'b0,x329 }<<<3'd1 )+$signed( { 3'b0,x330 }<<<3'd2 )+$signed( { 3'b0,x331 }<<<3'd2 )+$signed( -{ 3'b0,x332 }<<<3'd2)+$signed( { 4'b0,x333 }<<<3'd3 )+$signed( { 2'b0,x334 } <<<3'd1 )+$signed( { 3'b0,x335 }<<<3'd2 )+$signed( { 3'b0,x336 }<<<3'd2 )+$signed( { 2'b0,x337 } <<<3'd1 )+$signed( -{ 1'b0,x338 } )+$signed( { 2'b0,x340 } <<<3'd1 )+$signed( { 1'b0,x341 }  )+$signed( -{ 2'b0,x342 }<<<3'd1 )+$signed( -{ 1'b0,x343 } )+$signed( -{ 1'b0,x345 } )+$signed( { 2'b0,x346 } <<<3'd1 )+$signed( { 2'b0,x347 } <<<3'd1 )+$signed( -{ 3'b0,x349 }<<<3'd2)+$signed( { 1'b0,x350 }  )+$signed( -{ 1'b0,x351 } )+$signed( -{ 1'b0,x352 } )+$signed( { 2'b0,x353 } <<<3'd1 )+$signed( -{ 2'b0,x355 }<<<3'd1 )+$signed( -{ 1'b0,x356 } )+$signed( -{ 3'b0,x357 }<<<3'd2)+$signed( { 2'b0,x358 } <<<3'd1 )+$signed( -{ 1'b0,x359 } )+$signed( { 2'b0,x360 } <<<3'd1 )+$signed( { 2'b0,x361 } <<<3'd1 )+$signed( { 3'b0,x362 }<<<3'd2 )+$signed( -{ 1'b0,x365 } )+$signed( -{ 1'b0,x366 } )+$signed( -{ 1'b0,x368 } )+$signed( -{ 1'b0,x370 } )+$signed( { 4'b0,x371 }<<<3'd3 )+$signed( { 1'b0,x372 }  )+$signed( { 2'b0,x373 } <<<3'd1 )+$signed( -{ 2'b0,x374 }<<<3'd1 )+$signed( -{ 2'b0,x375 }<<<3'd1 )+$signed( { 1'b0,x376 }  )+$signed( -{ 2'b0,x377 }<<<3'd1 )+$signed( -{ 2'b0,x378 }<<<3'd1 )+$signed( -{ 2'b0,x379 }<<<3'd1 )+$signed( { 1'b0,x380 }  )+$signed( { 1'b0,x381 }  )+$signed( { 2'b0,x382 } <<<3'd1 )+$signed( { 3'b0,x383 }<<<3'd2 )+$signed( { 1'b0,x384 }  )+$signed( { 4'b0,x385 }<<<3'd3 )+$signed( { 1'b0,x386 }  )+$signed( { 2'b0,x387 } <<<3'd1 )+$signed( { 2'b0,x388 } <<<3'd1 )+$signed( -{ 2'b0,x389 }<<<3'd1 )+$signed( { 3'b0,x390 }<<<3'd2 )+$signed( -{ 3'b0,x391 }<<<3'd2)+$signed( -{ 3'b0,x392 }<<<3'd2)+$signed( { 3'b0,x393 }<<<3'd2 )+$signed( -{ 3'b0,x394 }<<<3'd2)+$signed( { 1'b0,x395 }  )+$signed( -{ 2'b0,x396 }<<<3'd1 )+$signed( -{ 3'b0,x397 }<<<3'd2)+$signed( { 1'b0,x398 }  )+$signed( { 1'b0,x399 }  )+$signed( { 4'b0,x400 }<<<3'd3 )+$signed( -{ 3'b0,x401 }<<<3'd2)+$signed( { 2'b0,x402 } <<<3'd1 )+$signed( -{ 4'b0, x403 }<<<3'd3 )+$signed( { 1'b0,x404 }  )+$signed( { 1'b0,x405 }  )+$signed( -{ 1'b0,x406 } )+$signed( { 3'b0,x407 }<<<3'd2 )+$signed( -{ 1'b0,x409 } )+$signed( -{ 1'b0,x410 } )+$signed( -{ 1'b0,x412 } )+$signed( { 1'b0,x413 }  )+$signed( -{ 4'b0, x414 }<<<3'd3 )+$signed( { 3'b0,x415 }<<<3'd2 )+$signed( { 3'b0,x416 }<<<3'd2 )+$signed( -{ 2'b0,x417 }<<<3'd1 )+$signed( { 1'b0,x418 }  )+$signed( { 1'b0,x419 }  )+$signed( { 3'b0,x420 }<<<3'd2 )+$signed( -{ 2'b0,x421 }<<<3'd1 )+$signed( -{ 3'b0,x422 }<<<3'd2)+$signed( { 1'b0,x423 }  )+$signed( { 1'b0,x424 }  )+$signed( -{ 1'b0,x425 } )+$signed( { 3'b0,x426 }<<<3'd2 )+$signed( -{ 3'b0,x427 }<<<3'd2)+$signed( { 2'b0,x428 } <<<3'd1 )+$signed( -{ 2'b0,x429 }<<<3'd1 )+$signed( { 2'b0,x430 } <<<3'd1 )+$signed( -{ 1'b0,x431 } )+$signed( -{ 2'b0,x432 }<<<3'd1 )+$signed( -{ 1'b0,x433 } )+$signed( -{ 2'b0,x434 }<<<3'd1 )+$signed( -{ 4'b0, x435 }<<<3'd3 )+$signed( -{ 1'b0,x436 } )+$signed( { 2'b0,x437 } <<<3'd1 )+$signed( { 1'b0,x438 }  )+$signed( { 3'b0,x439 }<<<3'd2 )+$signed( { 2'b0,x440 } <<<3'd1 )+$signed( { 1'b0,x441 }  )+$signed( -{ 3'b0,x442 }<<<3'd2)+$signed( { 3'b0,x443 }<<<3'd2 )+$signed( -{ 3'b0,x444 }<<<3'd2)+$signed( -{ 1'b0,x445 } )+$signed( -{ 3'b0,x446 }<<<3'd2)+$signed( { 3'b0,x447 }<<<3'd2 )+$signed( { 2'b0,x448 } <<<3'd1 )+$signed( -{ 3'b0,x449 }<<<3'd2)+$signed( -{ 2'b0,x450 }<<<3'd1 )+$signed( { 1'b0,x451 }  )+$signed( { 2'b0,x452 } <<<3'd1 )+$signed( -{ 2'b0,x454 }<<<3'd1 )+$signed( { 3'b0,x455 }<<<3'd2 )+$signed( { 1'b0,x456 }  )+$signed( -{ 2'b0,x457 }<<<3'd1 )+$signed( -{ 1'b0,x458 } )+$signed( -{ 3'b0,x459 }<<<3'd2)+$signed( { 4'b0,x460 }<<<3'd3 )+$signed( { 2'b0,x461 } <<<3'd1 )+$signed( { 2'b0,x462 } <<<3'd1 )+$signed( -{ 2'b0,x464 }<<<3'd1 )+$signed( -{ 3'b0,x465 }<<<3'd2)+$signed( -{ 3'b0,x467 }<<<3'd2)+$signed( { 3'b0,x468 }<<<3'd2 )+$signed( -{ 2'b0,x469 }<<<3'd1 )+$signed( { 3'b0,x470 }<<<3'd2 )+$signed( -{ 3'b0,x472 }<<<3'd2)+$signed( { 2'b0,x473 } <<<3'd1 )+$signed( -{ 2'b0,x474 }<<<3'd1 )+$signed( { 2'b0,x475 } <<<3'd1 )+$signed( { 2'b0,x477 } <<<3'd1 )+$signed( -{ 1'b0,x478 } )+$signed( { 2'b0,x479 } <<<3'd1 )+$signed( -{ 1'b0,x480 } )+$signed( { 2'b0,x481 } <<<3'd1 )+$signed( { 1'b0,x482 }  )+$signed( { 3'b0,x483 }<<<3'd2 )+$signed( { 1'b0,x484 }  )+$signed( -{ 1'b0,x485 } )+$signed( -{ 3'b0,x486 }<<<3'd2)+$signed( -{ 3'b0,x487 }<<<3'd2)+$signed( -{ 4'b0, x488 }<<<3'd3 )+$signed( -{ 2'b0,x489 }<<<3'd1 )+$signed( -{ 1'b0,x490 } )+$signed( -{ 3'b0,x491 }<<<3'd2)+$signed( { 3'b0,x492 }<<<3'd2 )+$signed( -{ 3'b0,x493 }<<<3'd2)+$signed( -{ 2'b0,x494 }<<<3'd1 )+$signed( -{ 2'b0,x495 }<<<3'd1 )+$signed(13'd16);
assign y7=temp_y[7][13] ==1'b1 ? 6'd0 :  
    temp_y[7][10] ==1'b1 ? 6'd63 : 
    temp_y[7][3]==1'b1 ? temp_y[7][9:4]+1'b1 : temp_y[7][9:4];
assign temp_y[8] = 
+$signed( -{ 2'b0,x0 }<<<3'd1 )+$signed( -{ 5'b0,x1 }<<<3'd4 )+$signed( { 3'b0,x2 }<<<3'd2 )+$signed( { 3'b0,x3 }<<<3'd2 )+$signed( { 4'b0,x4 }<<<3'd3 )+$signed( { 1'b0,x5 }  )+$signed( -{ 1'b0,x6 } )+$signed( -{ 5'b0,x8 }<<<3'd4 )+$signed( { 1'b0,x9 }  )+$signed( -{ 1'b0,x10 } )+$signed( -{ 3'b0,x11 }<<<3'd2)+$signed( { 2'b0,x12 } <<<3'd1 )+$signed( { 3'b0,x13 }<<<3'd2 )+$signed( -{ 3'b0,x14 }<<<3'd2)+$signed( { 3'b0,x15 }<<<3'd2 )+$signed( { 3'b0,x16 }<<<3'd2 )+$signed( -{ 2'b0,x17 }<<<3'd1 )+$signed( -{ 3'b0,x18 }<<<3'd2)+$signed( -{ 5'b0,x19 }<<<3'd4 )+$signed( { 3'b0,x20 }<<<3'd2 )+$signed( { 3'b0,x21 }<<<3'd2 )+$signed( { 3'b0,x22 }<<<3'd2 )+$signed( { 2'b0,x24 } <<<3'd1 )+$signed( { 2'b0,x25 } <<<3'd1 )+$signed( -{ 1'b0,x26 } )+$signed( { 1'b0,x27 }  )+$signed( -{ 3'b0,x28 }<<<3'd2)+$signed( -{ 3'b0,x29 }<<<3'd2)+$signed( { 1'b0,x30 }  )+$signed( { 2'b0,x31 } <<<3'd1 )+$signed( -{ 3'b0,x32 }<<<3'd2)+$signed( { 2'b0,x33 } <<<3'd1 )+$signed( -{ 1'b0,x34 } )+$signed( { 1'b0,x35 }  )+$signed( -{ 4'b0, x37 }<<<3'd3 )+$signed( { 3'b0,x38 }<<<3'd2 )+$signed( { 3'b0,x40 }<<<3'd2 )+$signed( { 2'b0,x42 } <<<3'd1 )+$signed( { 3'b0,x43 }<<<3'd2 )+$signed( -{ 4'b0, x44 }<<<3'd3 )+$signed( { 4'b0,x45 }<<<3'd3 )+$signed( -{ 3'b0,x46 }<<<3'd2)+$signed( -{ 3'b0,x47 }<<<3'd2)+$signed( -{ 3'b0,x48 }<<<3'd2)+$signed( { 1'b0,x49 }  )+$signed( -{ 2'b0,x50 }<<<3'd1 )+$signed( -{ 3'b0,x51 }<<<3'd2)+$signed( { 3'b0,x52 }<<<3'd2 )+$signed( { 3'b0,x53 }<<<3'd2 )+$signed( { 3'b0,x54 }<<<3'd2 )+$signed( -{ 4'b0, x55 }<<<3'd3 )+$signed( -{ 1'b0,x56 } )+$signed( { 1'b0,x57 }  )+$signed( { 2'b0,x59 } <<<3'd1 )+$signed( -{ 1'b0,x60 } )+$signed( { 2'b0,x61 } <<<3'd1 )+$signed( -{ 4'b0, x62 }<<<3'd3 )+$signed( { 3'b0,x63 }<<<3'd2 )+$signed( -{ 2'b0,x65 }<<<3'd1 )+$signed( { 3'b0,x66 }<<<3'd2 )+$signed( { 2'b0,x67 } <<<3'd1 )+$signed( { 3'b0,x69 }<<<3'd2 )+$signed( { 4'b0,x70 }<<<3'd3 )+$signed( { 3'b0,x71 }<<<3'd2 )+$signed( { 1'b0,x72 }  )+$signed( -{ 3'b0,x73 }<<<3'd2)+$signed( -{ 1'b0,x74 } )+$signed( -{ 3'b0,x75 }<<<3'd2)+$signed( { 3'b0,x76 }<<<3'd2 )+$signed( -{ 3'b0,x77 }<<<3'd2)+$signed( { 2'b0,x78 } <<<3'd1 )+$signed( { 3'b0,x79 }<<<3'd2 )+$signed( -{ 3'b0,x80 }<<<3'd2)+$signed( -{ 1'b0,x81 } )+$signed( { 1'b0,x82 }  )+$signed( -{ 2'b0,x83 }<<<3'd1 )+$signed( { 4'b0,x84 }<<<3'd3 )+$signed( { 3'b0,x85 }<<<3'd2 )+$signed( { 3'b0,x86 }<<<3'd2 )+$signed( { 1'b0,x88 }  )+$signed( { 3'b0,x89 }<<<3'd2 )+$signed( { 1'b0,x90 }  )+$signed( -{ 2'b0,x91 }<<<3'd1 )+$signed( { 3'b0,x93 }<<<3'd2 )+$signed( { 3'b0,x94 }<<<3'd2 )+$signed( -{ 2'b0,x95 }<<<3'd1 )+$signed( -{ 1'b0,x96 } )+$signed( -{ 2'b0,x97 }<<<3'd1 )+$signed( -{ 3'b0,x98 }<<<3'd2)+$signed( { 2'b0,x99 } <<<3'd1 )+$signed( -{ 3'b0,x100 }<<<3'd2)+$signed( { 1'b0,x101 }  )+$signed( { 2'b0,x102 } <<<3'd1 )+$signed( -{ 3'b0,x103 }<<<3'd2)+$signed( { 1'b0,x104 }  )+$signed( -{ 2'b0,x105 }<<<3'd1 )+$signed( -{ 3'b0,x106 }<<<3'd2)+$signed( -{ 2'b0,x107 }<<<3'd1 )+$signed( -{ 2'b0,x108 }<<<3'd1 )+$signed( -{ 3'b0,x109 }<<<3'd2)+$signed( { 3'b0,x111 }<<<3'd2 )+$signed( { 1'b0,x112 }  )+$signed( -{ 1'b0,x113 } )+$signed( -{ 1'b0,x114 } )+$signed( { 3'b0,x115 }<<<3'd2 )+$signed( -{ 5'b0,x116 }<<<3'd4 )+$signed( -{ 3'b0,x117 }<<<3'd2)+$signed( -{ 3'b0,x118 }<<<3'd2)+$signed( -{ 2'b0,x119 }<<<3'd1 )+$signed( -{ 3'b0,x121 }<<<3'd2)+$signed( -{ 3'b0,x122 }<<<3'd2)+$signed( { 2'b0,x123 } <<<3'd1 )+$signed( { 3'b0,x124 }<<<3'd2 )+$signed( -{ 3'b0,x125 }<<<3'd2)+$signed( { 3'b0,x126 }<<<3'd2 )+$signed( -{ 3'b0,x127 }<<<3'd2)+$signed( { 3'b0,x128 }<<<3'd2 )+$signed( -{ 3'b0,x129 }<<<3'd2)+$signed( -{ 2'b0,x130 }<<<3'd1 )+$signed( { 1'b0,x131 }  )+$signed( { 2'b0,x132 } <<<3'd1 )+$signed( -{ 2'b0,x133 }<<<3'd1 )+$signed( -{ 4'b0, x134 }<<<3'd3 )+$signed( -{ 2'b0,x136 }<<<3'd1 )+$signed( { 1'b0,x138 }  )+$signed( -{ 2'b0,x139 }<<<3'd1 )+$signed( -{ 2'b0,x140 }<<<3'd1 )+$signed( { 1'b0,x141 }  )+$signed( { 2'b0,x142 } <<<3'd1 )+$signed( { 2'b0,x143 } <<<3'd1 )+$signed( { 3'b0,x144 }<<<3'd2 )+$signed( -{ 3'b0,x145 }<<<3'd2)+$signed( -{ 1'b0,x146 } )+$signed( -{ 4'b0, x147 }<<<3'd3 )+$signed( -{ 3'b0,x149 }<<<3'd2)+$signed( -{ 1'b0,x150 } )+$signed( { 2'b0,x151 } <<<3'd1 )+$signed( -{ 2'b0,x152 }<<<3'd1 )+$signed( -{ 3'b0,x153 }<<<3'd2)+$signed( -{ 3'b0,x154 }<<<3'd2)+$signed( { 3'b0,x155 }<<<3'd2 )+$signed( -{ 3'b0,x156 }<<<3'd2)+$signed( -{ 2'b0,x157 }<<<3'd1 )+$signed( { 3'b0,x158 }<<<3'd2 )+$signed( -{ 1'b0,x159 } )+$signed( -{ 3'b0,x160 }<<<3'd2)+$signed( -{ 3'b0,x161 }<<<3'd2)+$signed( { 3'b0,x162 }<<<3'd2 )+$signed( { 3'b0,x163 }<<<3'd2 )+$signed( { 2'b0,x164 } <<<3'd1 )+$signed( { 3'b0,x165 }<<<3'd2 )+$signed( -{ 3'b0,x167 }<<<3'd2)+$signed( -{ 1'b0,x168 } )+$signed( -{ 1'b0,x169 } )+$signed( -{ 1'b0,x170 } )+$signed( -{ 3'b0,x171 }<<<3'd2)+$signed( { 2'b0,x173 } <<<3'd1 )+$signed( -{ 1'b0,x174 } )+$signed( -{ 3'b0,x176 }<<<3'd2)+$signed( -{ 1'b0,x177 } )+$signed( { 2'b0,x178 } <<<3'd1 )+$signed( -{ 2'b0,x179 }<<<3'd1 )+$signed( { 2'b0,x180 } <<<3'd1 )+$signed( { 3'b0,x181 }<<<3'd2 )+$signed( -{ 1'b0,x182 } )+$signed( { 1'b0,x183 }  )+$signed( { 2'b0,x185 } <<<3'd1 )+$signed( { 2'b0,x188 } <<<3'd1 )+$signed( -{ 3'b0,x189 }<<<3'd2)+$signed( { 3'b0,x190 }<<<3'd2 )+$signed( { 3'b0,x191 }<<<3'd2 )+$signed( { 1'b0,x192 }  )+$signed( { 3'b0,x193 }<<<3'd2 )+$signed( { 1'b0,x194 }  )+$signed( -{ 2'b0,x196 }<<<3'd1 )+$signed( { 2'b0,x197 } <<<3'd1 )+$signed( { 3'b0,x199 }<<<3'd2 )+$signed( -{ 3'b0,x200 }<<<3'd2)+$signed( { 2'b0,x201 } <<<3'd1 )+$signed( -{ 3'b0,x202 }<<<3'd2)+$signed( -{ 2'b0,x203 }<<<3'd1 )+$signed( -{ 1'b0,x204 } )+$signed( { 1'b0,x205 }  )+$signed( -{ 1'b0,x206 } )+$signed( -{ 3'b0,x207 }<<<3'd2)+$signed( { 3'b0,x208 }<<<3'd2 )+$signed( { 1'b0,x209 }  )+$signed( { 1'b0,x210 }  )+$signed( { 3'b0,x211 }<<<3'd2 )+$signed( { 2'b0,x212 } <<<3'd1 )+$signed( -{ 1'b0,x213 } )+$signed( { 2'b0,x214 } <<<3'd1 )+$signed( -{ 2'b0,x215 }<<<3'd1 )+$signed( { 2'b0,x216 } <<<3'd1 )+$signed( -{ 2'b0,x217 }<<<3'd1 )+$signed( -{ 2'b0,x218 }<<<3'd1 )+$signed( -{ 2'b0,x219 }<<<3'd1 )+$signed( { 1'b0,x220 }  )+$signed( -{ 3'b0,x221 }<<<3'd2)+$signed( { 2'b0,x222 } <<<3'd1 )+$signed( -{ 3'b0,x223 }<<<3'd2)+$signed( -{ 4'b0, x224 }<<<3'd3 )+$signed( { 2'b0,x225 } <<<3'd1 )+$signed( -{ 2'b0,x226 }<<<3'd1 )+$signed( -{ 2'b0,x227 }<<<3'd1 )+$signed( { 2'b0,x228 } <<<3'd1 )+$signed( -{ 3'b0,x231 }<<<3'd2)+$signed( { 1'b0,x232 }  )+$signed( -{ 1'b0,x233 } )+$signed( -{ 1'b0,x234 } )+$signed( { 3'b0,x235 }<<<3'd2 )+$signed( -{ 2'b0,x236 }<<<3'd1 )+$signed( { 3'b0,x237 }<<<3'd2 )+$signed( { 2'b0,x238 } <<<3'd1 )+$signed( -{ 2'b0,x239 }<<<3'd1 )+$signed( { 1'b0,x240 }  )+$signed( { 3'b0,x241 }<<<3'd2 )+$signed( -{ 4'b0, x242 }<<<3'd3 )+$signed( -{ 4'b0, x243 }<<<3'd3 )+$signed( -{ 3'b0,x244 }<<<3'd2)+$signed( { 3'b0,x245 }<<<3'd2 )+$signed( -{ 2'b0,x246 }<<<3'd1 )+$signed( -{ 2'b0,x247 }<<<3'd1 )+$signed( { 1'b0,x248 }  )+$signed( -{ 1'b0,x249 } )+$signed( { 2'b0,x250 } <<<3'd1 )+$signed( -{ 2'b0,x251 }<<<3'd1 )+$signed( { 2'b0,x252 } <<<3'd1 )+$signed( { 4'b0,x253 }<<<3'd3 )+$signed( { 2'b0,x254 } <<<3'd1 )+$signed( { 3'b0,x255 }<<<3'd2 )+$signed( -{ 3'b0,x257 }<<<3'd2)+$signed( { 2'b0,x258 } <<<3'd1 )+$signed( { 1'b0,x259 }  )+$signed( -{ 2'b0,x260 }<<<3'd1 )+$signed( -{ 5'b0,x261 }<<<3'd4 )+$signed( -{ 3'b0,x262 }<<<3'd2)+$signed( { 1'b0,x263 }  )+$signed( -{ 3'b0,x264 }<<<3'd2)+$signed( -{ 3'b0,x265 }<<<3'd2)+$signed( -{ 1'b0,x266 } )+$signed( -{ 1'b0,x267 } )+$signed( { 2'b0,x268 } <<<3'd1 )+$signed( { 2'b0,x269 } <<<3'd1 )+$signed( { 2'b0,x270 } <<<3'd1 )+$signed( { 2'b0,x271 } <<<3'd1 )+$signed( { 3'b0,x273 }<<<3'd2 )+$signed( { 3'b0,x274 }<<<3'd2 )+$signed( -{ 2'b0,x275 }<<<3'd1 )+$signed( { 2'b0,x276 } <<<3'd1 )+$signed( { 2'b0,x277 } <<<3'd1 )+$signed( -{ 4'b0, x278 }<<<3'd3 )+$signed( -{ 4'b0, x279 }<<<3'd3 )+$signed( { 3'b0,x280 }<<<3'd2 )+$signed( { 1'b0,x281 }  )+$signed( -{ 3'b0,x282 }<<<3'd2)+$signed( -{ 1'b0,x283 } )+$signed( -{ 2'b0,x285 }<<<3'd1 )+$signed( -{ 2'b0,x286 }<<<3'd1 )+$signed( { 2'b0,x287 } <<<3'd1 )+$signed( { 2'b0,x288 } <<<3'd1 )+$signed( { 3'b0,x289 }<<<3'd2 )+$signed( { 3'b0,x290 }<<<3'd2 )+$signed( { 4'b0,x291 }<<<3'd3 )+$signed( { 4'b0,x292 }<<<3'd3 )+$signed( -{ 2'b0,x293 }<<<3'd1 )+$signed( { 2'b0,x294 } <<<3'd1 )+$signed( -{ 3'b0,x295 }<<<3'd2)+$signed( -{ 4'b0, x296 }<<<3'd3 )+$signed( -{ 1'b0,x297 } )+$signed( -{ 2'b0,x298 }<<<3'd1 )+$signed( -{ 1'b0,x299 } )+$signed( { 3'b0,x300 }<<<3'd2 )+$signed( -{ 1'b0,x301 } )+$signed( { 2'b0,x302 } <<<3'd1 )+$signed( -{ 1'b0,x303 } )+$signed( { 3'b0,x304 }<<<3'd2 )+$signed( { 1'b0,x305 }  )+$signed( -{ 3'b0,x306 }<<<3'd2)+$signed( -{ 1'b0,x307 } )+$signed( -{ 3'b0,x308 }<<<3'd2)+$signed( { 2'b0,x309 } <<<3'd1 )+$signed( -{ 4'b0, x310 }<<<3'd3 )+$signed( { 3'b0,x311 }<<<3'd2 )+$signed( { 2'b0,x312 } <<<3'd1 )+$signed( { 3'b0,x313 }<<<3'd2 )+$signed( { 2'b0,x314 } <<<3'd1 )+$signed( { 3'b0,x315 }<<<3'd2 )+$signed( { 2'b0,x316 } <<<3'd1 )+$signed( -{ 2'b0,x317 }<<<3'd1 )+$signed( -{ 2'b0,x318 }<<<3'd1 )+$signed( -{ 2'b0,x319 }<<<3'd1 )+$signed( { 4'b0,x320 }<<<3'd3 )+$signed( { 1'b0,x321 }  )+$signed( -{ 3'b0,x323 }<<<3'd2)+$signed( { 1'b0,x324 }  )+$signed( -{ 3'b0,x325 }<<<3'd2)+$signed( { 2'b0,x326 } <<<3'd1 )+$signed( { 2'b0,x328 } <<<3'd1 )+$signed( { 3'b0,x329 }<<<3'd2 )+$signed( -{ 1'b0,x330 } )+$signed( -{ 2'b0,x331 }<<<3'd1 )+$signed( { 3'b0,x332 }<<<3'd2 )+$signed( { 1'b0,x334 }  )+$signed( { 3'b0,x335 }<<<3'd2 )+$signed( -{ 2'b0,x336 }<<<3'd1 )+$signed( { 4'b0,x337 }<<<3'd3 )+$signed( { 2'b0,x338 } <<<3'd1 )+$signed( { 4'b0,x339 }<<<3'd3 )+$signed( -{ 1'b0,x341 } )+$signed( { 3'b0,x342 }<<<3'd2 )+$signed( { 1'b0,x343 }  )+$signed( -{ 4'b0, x344 }<<<3'd3 )+$signed( -{ 3'b0,x345 }<<<3'd2)+$signed( -{ 2'b0,x346 }<<<3'd1 )+$signed( -{ 3'b0,x347 }<<<3'd2)+$signed( -{ 3'b0,x348 }<<<3'd2)+$signed( -{ 1'b0,x349 } )+$signed( { 2'b0,x352 } <<<3'd1 )+$signed( -{ 4'b0, x356 }<<<3'd3 )+$signed( -{ 1'b0,x357 } )+$signed( -{ 2'b0,x358 }<<<3'd1 )+$signed( -{ 1'b0,x360 } )+$signed( { 2'b0,x361 } <<<3'd1 )+$signed( -{ 5'b0,x362 }<<<3'd4 )+$signed( { 3'b0,x364 }<<<3'd2 )+$signed( { 4'b0,x365 }<<<3'd3 )+$signed( -{ 3'b0,x366 }<<<3'd2)+$signed( { 1'b0,x367 }  )+$signed( -{ 1'b0,x368 } )+$signed( -{ 3'b0,x369 }<<<3'd2)+$signed( { 1'b0,x370 }  )+$signed( -{ 3'b0,x371 }<<<3'd2)+$signed( { 2'b0,x372 } <<<3'd1 )+$signed( -{ 1'b0,x374 } )+$signed( -{ 5'b0,x375 }<<<3'd4 )+$signed( -{ 5'b0,x377 }<<<3'd4 )+$signed( -{ 1'b0,x380 } )+$signed( { 2'b0,x381 } <<<3'd1 )+$signed( -{ 1'b0,x382 } )+$signed( -{ 1'b0,x383 } )+$signed( { 3'b0,x385 }<<<3'd2 )+$signed( { 2'b0,x386 } <<<3'd1 )+$signed( { 3'b0,x387 }<<<3'd2 )+$signed( -{ 4'b0, x388 }<<<3'd3 )+$signed( { 2'b0,x389 } <<<3'd1 )+$signed( -{ 1'b0,x390 } )+$signed( { 2'b0,x391 } <<<3'd1 )+$signed( { 3'b0,x393 }<<<3'd2 )+$signed( { 2'b0,x394 } <<<3'd1 )+$signed( -{ 2'b0,x396 }<<<3'd1 )+$signed( { 1'b0,x397 }  )+$signed( { 2'b0,x398 } <<<3'd1 )+$signed( { 2'b0,x400 } <<<3'd1 )+$signed( -{ 3'b0,x402 }<<<3'd2)+$signed( { 3'b0,x403 }<<<3'd2 )+$signed( { 2'b0,x406 } <<<3'd1 )+$signed( { 3'b0,x407 }<<<3'd2 )+$signed( { 1'b0,x409 }  )+$signed( { 2'b0,x410 } <<<3'd1 )+$signed( { 2'b0,x411 } <<<3'd1 )+$signed( -{ 1'b0,x412 } )+$signed( -{ 3'b0,x414 }<<<3'd2)+$signed( -{ 2'b0,x415 }<<<3'd1 )+$signed( { 2'b0,x416 } <<<3'd1 )+$signed( { 2'b0,x418 } <<<3'd1 )+$signed( { 1'b0,x419 }  )+$signed( -{ 3'b0,x420 }<<<3'd2)+$signed( { 2'b0,x421 } <<<3'd1 )+$signed( -{ 1'b0,x422 } )+$signed( { 2'b0,x423 } <<<3'd1 )+$signed( -{ 1'b0,x424 } )+$signed( -{ 1'b0,x425 } )+$signed( { 1'b0,x426 }  )+$signed( -{ 5'b0,x427 }<<<3'd4 )+$signed( -{ 1'b0,x428 } )+$signed( { 2'b0,x429 } <<<3'd1 )+$signed( { 2'b0,x430 } <<<3'd1 )+$signed( -{ 2'b0,x431 }<<<3'd1 )+$signed( -{ 2'b0,x432 }<<<3'd1 )+$signed( { 1'b0,x433 }  )+$signed( { 1'b0,x434 }  )+$signed( -{ 1'b0,x435 } )+$signed( { 1'b0,x436 }  )+$signed( { 3'b0,x437 }<<<3'd2 )+$signed( -{ 2'b0,x438 }<<<3'd1 )+$signed( -{ 2'b0,x439 }<<<3'd1 )+$signed( -{ 3'b0,x440 }<<<3'd2)+$signed( { 2'b0,x442 } <<<3'd1 )+$signed( { 3'b0,x443 }<<<3'd2 )+$signed( { 1'b0,x444 }  )+$signed( { 1'b0,x445 }  )+$signed( { 3'b0,x446 }<<<3'd2 )+$signed( -{ 2'b0,x447 }<<<3'd1 )+$signed( -{ 1'b0,x448 } )+$signed( -{ 1'b0,x449 } )+$signed( -{ 1'b0,x451 } )+$signed( -{ 1'b0,x452 } )+$signed( -{ 3'b0,x453 }<<<3'd2)+$signed( -{ 2'b0,x454 }<<<3'd1 )+$signed( { 3'b0,x455 }<<<3'd2 )+$signed( { 3'b0,x457 }<<<3'd2 )+$signed( { 2'b0,x458 } <<<3'd1 )+$signed( { 3'b0,x459 }<<<3'd2 )+$signed( { 3'b0,x460 }<<<3'd2 )+$signed( -{ 1'b0,x462 } )+$signed( -{ 1'b0,x463 } )+$signed( { 1'b0,x464 }  )+$signed( -{ 2'b0,x466 }<<<3'd1 )+$signed( { 2'b0,x467 } <<<3'd1 )+$signed( { 3'b0,x468 }<<<3'd2 )+$signed( { 3'b0,x469 }<<<3'd2 )+$signed( { 2'b0,x470 } <<<3'd1 )+$signed( { 2'b0,x471 } <<<3'd1 )+$signed( { 4'b0,x472 }<<<3'd3 )+$signed( { 2'b0,x473 } <<<3'd1 )+$signed( { 2'b0,x474 } <<<3'd1 )+$signed( -{ 2'b0,x475 }<<<3'd1 )+$signed( { 1'b0,x476 }  )+$signed( { 2'b0,x477 } <<<3'd1 )+$signed( -{ 2'b0,x478 }<<<3'd1 )+$signed( -{ 3'b0,x479 }<<<3'd2)+$signed( -{ 3'b0,x480 }<<<3'd2)+$signed( { 1'b0,x481 }  )+$signed( { 1'b0,x482 }  )+$signed( { 2'b0,x483 } <<<3'd1 )+$signed( { 3'b0,x484 }<<<3'd2 )+$signed( { 2'b0,x485 } <<<3'd1 )+$signed( -{ 1'b0,x486 } )+$signed( -{ 1'b0,x487 } )+$signed( { 1'b0,x488 }  )+$signed( { 1'b0,x489 }  )+$signed( { 3'b0,x490 }<<<3'd2 )+$signed( -{ 4'b0, x491 }<<<3'd3 )+$signed( -{ 4'b0, x492 }<<<3'd3 )+$signed( { 1'b0,x493 }  )+$signed( -{ 1'b0,x494 } )+$signed( { 4'b0,x495 }<<<3'd3 )+$signed(13'd24);
assign y8=temp_y[8][13] ==1'b1 ? 6'd0 :  
    temp_y[8][10] ==1'b1 ? 6'd63 : 
    temp_y[8][3]==1'b1 ? temp_y[8][9:4]+1'b1 : temp_y[8][9:4];
assign temp_y[9] = 
+$signed( { 3'b0,x0 }<<<3'd2 )+$signed( { 1'b0,x1 }  )+$signed( -{ 1'b0,x3 } )+$signed( -{ 2'b0,x4 }<<<3'd1 )+$signed( -{ 2'b0,x5 }<<<3'd1 )+$signed( { 1'b0,x6 }  )+$signed( { 4'b0,x7 }<<<3'd3 )+$signed( { 4'b0,x8 }<<<3'd3 )+$signed( { 1'b0,x11 }  )+$signed( -{ 2'b0,x12 }<<<3'd1 )+$signed( { 1'b0,x13 }  )+$signed( -{ 2'b0,x14 }<<<3'd1 )+$signed( { 2'b0,x15 } <<<3'd1 )+$signed( -{ 4'b0, x16 }<<<3'd3 )+$signed( -{ 2'b0,x17 }<<<3'd1 )+$signed( { 3'b0,x18 }<<<3'd2 )+$signed( -{ 1'b0,x19 } )+$signed( -{ 3'b0,x20 }<<<3'd2)+$signed( { 3'b0,x21 }<<<3'd2 )+$signed( -{ 3'b0,x22 }<<<3'd2)+$signed( -{ 1'b0,x24 } )+$signed( { 3'b0,x25 }<<<3'd2 )+$signed( { 3'b0,x26 }<<<3'd2 )+$signed( -{ 3'b0,x27 }<<<3'd2)+$signed( -{ 2'b0,x28 }<<<3'd1 )+$signed( { 1'b0,x29 }  )+$signed( -{ 2'b0,x30 }<<<3'd1 )+$signed( { 2'b0,x31 } <<<3'd1 )+$signed( { 5'b0,x32  }<<<3'd4 )+$signed( -{ 3'b0,x33 }<<<3'd2)+$signed( -{ 1'b0,x34 } )+$signed( { 1'b0,x35 }  )+$signed( -{ 2'b0,x37 }<<<3'd1 )+$signed( -{ 3'b0,x38 }<<<3'd2)+$signed( { 2'b0,x39 } <<<3'd1 )+$signed( -{ 3'b0,x40 }<<<3'd2)+$signed( { 1'b0,x41 }  )+$signed( { 2'b0,x42 } <<<3'd1 )+$signed( { 2'b0,x43 } <<<3'd1 )+$signed( { 3'b0,x44 }<<<3'd2 )+$signed( -{ 2'b0,x45 }<<<3'd1 )+$signed( -{ 1'b0,x47 } )+$signed( -{ 3'b0,x48 }<<<3'd2)+$signed( { 4'b0,x50 }<<<3'd3 )+$signed( -{ 4'b0, x51 }<<<3'd3 )+$signed( { 2'b0,x54 } <<<3'd1 )+$signed( -{ 2'b0,x55 }<<<3'd1 )+$signed( -{ 1'b0,x56 } )+$signed( { 1'b0,x57 }  )+$signed( -{ 2'b0,x58 }<<<3'd1 )+$signed( -{ 2'b0,x59 }<<<3'd1 )+$signed( -{ 1'b0,x60 } )+$signed( { 1'b0,x61 }  )+$signed( { 1'b0,x62 }  )+$signed( { 1'b0,x65 }  )+$signed( -{ 3'b0,x66 }<<<3'd2)+$signed( -{ 1'b0,x68 } )+$signed( -{ 2'b0,x69 }<<<3'd1 )+$signed( { 2'b0,x71 } <<<3'd1 )+$signed( { 1'b0,x72 }  )+$signed( { 2'b0,x73 } <<<3'd1 )+$signed( { 2'b0,x74 } <<<3'd1 )+$signed( -{ 1'b0,x75 } )+$signed( { 3'b0,x76 }<<<3'd2 )+$signed( { 2'b0,x77 } <<<3'd1 )+$signed( -{ 1'b0,x78 } )+$signed( -{ 2'b0,x81 }<<<3'd1 )+$signed( -{ 1'b0,x82 } )+$signed( { 1'b0,x83 }  )+$signed( -{ 3'b0,x84 }<<<3'd2)+$signed( -{ 3'b0,x86 }<<<3'd2)+$signed( { 2'b0,x87 } <<<3'd1 )+$signed( { 3'b0,x88 }<<<3'd2 )+$signed( { 2'b0,x90 } <<<3'd1 )+$signed( { 1'b0,x91 }  )+$signed( -{ 3'b0,x92 }<<<3'd2)+$signed( { 3'b0,x93 }<<<3'd2 )+$signed( { 2'b0,x94 } <<<3'd1 )+$signed( { 1'b0,x95 }  )+$signed( -{ 4'b0, x97 }<<<3'd3 )+$signed( -{ 2'b0,x98 }<<<3'd1 )+$signed( { 2'b0,x99 } <<<3'd1 )+$signed( { 2'b0,x100 } <<<3'd1 )+$signed( -{ 3'b0,x101 }<<<3'd2)+$signed( { 1'b0,x103 }  )+$signed( -{ 3'b0,x105 }<<<3'd2)+$signed( { 2'b0,x107 } <<<3'd1 )+$signed( { 3'b0,x108 }<<<3'd2 )+$signed( -{ 2'b0,x109 }<<<3'd1 )+$signed( { 2'b0,x110 } <<<3'd1 )+$signed( { 3'b0,x111 }<<<3'd2 )+$signed( -{ 3'b0,x112 }<<<3'd2)+$signed( { 1'b0,x113 }  )+$signed( { 2'b0,x114 } <<<3'd1 )+$signed( { 3'b0,x115 }<<<3'd2 )+$signed( -{ 2'b0,x116 }<<<3'd1 )+$signed( -{ 2'b0,x117 }<<<3'd1 )+$signed( { 3'b0,x118 }<<<3'd2 )+$signed( { 2'b0,x119 } <<<3'd1 )+$signed( -{ 1'b0,x120 } )+$signed( -{ 2'b0,x121 }<<<3'd1 )+$signed( -{ 2'b0,x123 }<<<3'd1 )+$signed( -{ 3'b0,x124 }<<<3'd2)+$signed( { 2'b0,x125 } <<<3'd1 )+$signed( -{ 3'b0,x126 }<<<3'd2)+$signed( -{ 2'b0,x127 }<<<3'd1 )+$signed( -{ 2'b0,x128 }<<<3'd1 )+$signed( { 1'b0,x129 }  )+$signed( { 3'b0,x133 }<<<3'd2 )+$signed( -{ 2'b0,x134 }<<<3'd1 )+$signed( { 3'b0,x135 }<<<3'd2 )+$signed( -{ 1'b0,x138 } )+$signed( { 2'b0,x139 } <<<3'd1 )+$signed( { 2'b0,x141 } <<<3'd1 )+$signed( -{ 3'b0,x142 }<<<3'd2)+$signed( { 2'b0,x143 } <<<3'd1 )+$signed( { 3'b0,x144 }<<<3'd2 )+$signed( -{ 2'b0,x145 }<<<3'd1 )+$signed( -{ 3'b0,x146 }<<<3'd2)+$signed( -{ 2'b0,x147 }<<<3'd1 )+$signed( -{ 3'b0,x148 }<<<3'd2)+$signed( { 1'b0,x149 }  )+$signed( { 1'b0,x150 }  )+$signed( -{ 3'b0,x151 }<<<3'd2)+$signed( { 1'b0,x152 }  )+$signed( { 1'b0,x153 }  )+$signed( -{ 2'b0,x154 }<<<3'd1 )+$signed( -{ 2'b0,x155 }<<<3'd1 )+$signed( { 2'b0,x157 } <<<3'd1 )+$signed( { 3'b0,x158 }<<<3'd2 )+$signed( { 2'b0,x159 } <<<3'd1 )+$signed( { 2'b0,x160 } <<<3'd1 )+$signed( -{ 1'b0,x162 } )+$signed( { 3'b0,x163 }<<<3'd2 )+$signed( -{ 3'b0,x164 }<<<3'd2)+$signed( -{ 2'b0,x165 }<<<3'd1 )+$signed( { 1'b0,x166 }  )+$signed( { 1'b0,x167 }  )+$signed( -{ 3'b0,x169 }<<<3'd2)+$signed( { 2'b0,x171 } <<<3'd1 )+$signed( { 1'b0,x172 }  )+$signed( { 3'b0,x173 }<<<3'd2 )+$signed( { 3'b0,x174 }<<<3'd2 )+$signed( -{ 1'b0,x175 } )+$signed( { 2'b0,x176 } <<<3'd1 )+$signed( -{ 1'b0,x177 } )+$signed( { 2'b0,x178 } <<<3'd1 )+$signed( -{ 4'b0, x180 }<<<3'd3 )+$signed( { 3'b0,x181 }<<<3'd2 )+$signed( -{ 3'b0,x182 }<<<3'd2)+$signed( -{ 2'b0,x183 }<<<3'd1 )+$signed( -{ 3'b0,x184 }<<<3'd2)+$signed( -{ 1'b0,x185 } )+$signed( -{ 2'b0,x186 }<<<3'd1 )+$signed( -{ 3'b0,x187 }<<<3'd2)+$signed( -{ 2'b0,x189 }<<<3'd1 )+$signed( { 1'b0,x190 }  )+$signed( -{ 2'b0,x191 }<<<3'd1 )+$signed( { 3'b0,x192 }<<<3'd2 )+$signed( { 1'b0,x193 }  )+$signed( { 2'b0,x194 } <<<3'd1 )+$signed( -{ 2'b0,x195 }<<<3'd1 )+$signed( { 3'b0,x196 }<<<3'd2 )+$signed( { 2'b0,x197 } <<<3'd1 )+$signed( -{ 1'b0,x199 } )+$signed( -{ 4'b0, x200 }<<<3'd3 )+$signed( -{ 1'b0,x201 } )+$signed( -{ 3'b0,x202 }<<<3'd2)+$signed( { 2'b0,x203 } <<<3'd1 )+$signed( -{ 3'b0,x205 }<<<3'd2)+$signed( -{ 1'b0,x206 } )+$signed( { 3'b0,x207 }<<<3'd2 )+$signed( { 1'b0,x210 }  )+$signed( { 2'b0,x211 } <<<3'd1 )+$signed( { 1'b0,x212 }  )+$signed( -{ 4'b0, x213 }<<<3'd3 )+$signed( { 2'b0,x214 } <<<3'd1 )+$signed( -{ 2'b0,x215 }<<<3'd1 )+$signed( -{ 3'b0,x216 }<<<3'd2)+$signed( -{ 4'b0, x217 }<<<3'd3 )+$signed( -{ 3'b0,x218 }<<<3'd2)+$signed( { 3'b0,x219 }<<<3'd2 )+$signed( { 2'b0,x220 } <<<3'd1 )+$signed( -{ 2'b0,x221 }<<<3'd1 )+$signed( { 2'b0,x222 } <<<3'd1 )+$signed( { 3'b0,x223 }<<<3'd2 )+$signed( { 3'b0,x224 }<<<3'd2 )+$signed( { 3'b0,x225 }<<<3'd2 )+$signed( -{ 3'b0,x226 }<<<3'd2)+$signed( -{ 2'b0,x227 }<<<3'd1 )+$signed( { 2'b0,x228 } <<<3'd1 )+$signed( { 3'b0,x229 }<<<3'd2 )+$signed( { 1'b0,x230 }  )+$signed( { 2'b0,x231 } <<<3'd1 )+$signed( { 2'b0,x232 } <<<3'd1 )+$signed( -{ 1'b0,x233 } )+$signed( -{ 2'b0,x234 }<<<3'd1 )+$signed( -{ 3'b0,x235 }<<<3'd2)+$signed( -{ 2'b0,x236 }<<<3'd1 )+$signed( { 2'b0,x237 } <<<3'd1 )+$signed( -{ 3'b0,x238 }<<<3'd2)+$signed( -{ 2'b0,x239 }<<<3'd1 )+$signed( { 2'b0,x240 } <<<3'd1 )+$signed( { 3'b0,x241 }<<<3'd2 )+$signed( { 2'b0,x242 } <<<3'd1 )+$signed( { 3'b0,x243 }<<<3'd2 )+$signed( -{ 4'b0, x244 }<<<3'd3 )+$signed( -{ 1'b0,x245 } )+$signed( { 2'b0,x246 } <<<3'd1 )+$signed( { 1'b0,x247 }  )+$signed( { 3'b0,x248 }<<<3'd2 )+$signed( -{ 3'b0,x249 }<<<3'd2)+$signed( { 3'b0,x250 }<<<3'd2 )+$signed( -{ 3'b0,x251 }<<<3'd2)+$signed( -{ 3'b0,x252 }<<<3'd2)+$signed( -{ 4'b0, x253 }<<<3'd3 )+$signed( { 1'b0,x254 }  )+$signed( -{ 3'b0,x255 }<<<3'd2)+$signed( -{ 3'b0,x256 }<<<3'd2)+$signed( -{ 1'b0,x257 } )+$signed( { 2'b0,x258 } <<<3'd1 )+$signed( { 1'b0,x259 }  )+$signed( { 3'b0,x260 }<<<3'd2 )+$signed( -{ 2'b0,x262 }<<<3'd1 )+$signed( -{ 3'b0,x264 }<<<3'd2)+$signed( { 2'b0,x265 } <<<3'd1 )+$signed( { 3'b0,x266 }<<<3'd2 )+$signed( -{ 4'b0, x267 }<<<3'd3 )+$signed( { 2'b0,x268 } <<<3'd1 )+$signed( -{ 2'b0,x269 }<<<3'd1 )+$signed( -{ 3'b0,x270 }<<<3'd2)+$signed( -{ 3'b0,x271 }<<<3'd2)+$signed( -{ 4'b0, x272 }<<<3'd3 )+$signed( -{ 1'b0,x273 } )+$signed( -{ 3'b0,x274 }<<<3'd2)+$signed( -{ 2'b0,x275 }<<<3'd1 )+$signed( { 2'b0,x276 } <<<3'd1 )+$signed( { 3'b0,x277 }<<<3'd2 )+$signed( { 3'b0,x278 }<<<3'd2 )+$signed( { 3'b0,x279 }<<<3'd2 )+$signed( -{ 4'b0, x280 }<<<3'd3 )+$signed( -{ 2'b0,x281 }<<<3'd1 )+$signed( { 1'b0,x282 }  )+$signed( { 3'b0,x284 }<<<3'd2 )+$signed( -{ 3'b0,x286 }<<<3'd2)+$signed( { 2'b0,x287 } <<<3'd1 )+$signed( { 2'b0,x288 } <<<3'd1 )+$signed( { 2'b0,x289 } <<<3'd1 )+$signed( { 3'b0,x290 }<<<3'd2 )+$signed( -{ 2'b0,x291 }<<<3'd1 )+$signed( -{ 3'b0,x293 }<<<3'd2)+$signed( -{ 4'b0, x294 }<<<3'd3 )+$signed( -{ 2'b0,x295 }<<<3'd1 )+$signed( { 3'b0,x296 }<<<3'd2 )+$signed( { 2'b0,x297 } <<<3'd1 )+$signed( -{ 2'b0,x298 }<<<3'd1 )+$signed( { 3'b0,x299 }<<<3'd2 )+$signed( { 2'b0,x301 } <<<3'd1 )+$signed( -{ 4'b0, x302 }<<<3'd3 )+$signed( { 3'b0,x303 }<<<3'd2 )+$signed( { 1'b0,x304 }  )+$signed( -{ 3'b0,x305 }<<<3'd2)+$signed( { 2'b0,x306 } <<<3'd1 )+$signed( -{ 4'b0, x307 }<<<3'd3 )+$signed( -{ 3'b0,x308 }<<<3'd2)+$signed( { 3'b0,x309 }<<<3'd2 )+$signed( -{ 2'b0,x310 }<<<3'd1 )+$signed( -{ 4'b0, x311 }<<<3'd3 )+$signed( { 3'b0,x312 }<<<3'd2 )+$signed( { 1'b0,x314 }  )+$signed( -{ 4'b0, x315 }<<<3'd3 )+$signed( { 3'b0,x316 }<<<3'd2 )+$signed( -{ 2'b0,x317 }<<<3'd1 )+$signed( -{ 1'b0,x318 } )+$signed( -{ 3'b0,x320 }<<<3'd2)+$signed( -{ 3'b0,x321 }<<<3'd2)+$signed( -{ 3'b0,x322 }<<<3'd2)+$signed( -{ 3'b0,x323 }<<<3'd2)+$signed( -{ 4'b0, x324 }<<<3'd3 )+$signed( { 1'b0,x325 }  )+$signed( -{ 3'b0,x328 }<<<3'd2)+$signed( { 3'b0,x329 }<<<3'd2 )+$signed( -{ 2'b0,x330 }<<<3'd1 )+$signed( -{ 3'b0,x332 }<<<3'd2)+$signed( -{ 2'b0,x333 }<<<3'd1 )+$signed( -{ 3'b0,x334 }<<<3'd2)+$signed( -{ 3'b0,x335 }<<<3'd2)+$signed( { 1'b0,x336 }  )+$signed( -{ 4'b0, x337 }<<<3'd3 )+$signed( { 1'b0,x338 }  )+$signed( -{ 3'b0,x339 }<<<3'd2)+$signed( { 1'b0,x340 }  )+$signed( -{ 2'b0,x341 }<<<3'd1 )+$signed( -{ 1'b0,x343 } )+$signed( { 3'b0,x344 }<<<3'd2 )+$signed( -{ 1'b0,x345 } )+$signed( { 2'b0,x346 } <<<3'd1 )+$signed( { 3'b0,x347 }<<<3'd2 )+$signed( { 1'b0,x348 }  )+$signed( { 1'b0,x349 }  )+$signed( { 3'b0,x350 }<<<3'd2 )+$signed( -{ 2'b0,x351 }<<<3'd1 )+$signed( -{ 3'b0,x352 }<<<3'd2)+$signed( { 2'b0,x353 } <<<3'd1 )+$signed( { 3'b0,x354 }<<<3'd2 )+$signed( { 3'b0,x355 }<<<3'd2 )+$signed( -{ 1'b0,x356 } )+$signed( { 3'b0,x357 }<<<3'd2 )+$signed( -{ 4'b0, x359 }<<<3'd3 )+$signed( { 2'b0,x360 } <<<3'd1 )+$signed( -{ 2'b0,x361 }<<<3'd1 )+$signed( { 4'b0,x362 }<<<3'd3 )+$signed( -{ 4'b0, x363 }<<<3'd3 )+$signed( { 3'b0,x364 }<<<3'd2 )+$signed( -{ 4'b0, x365 }<<<3'd3 )+$signed( { 3'b0,x366 }<<<3'd2 )+$signed( { 3'b0,x367 }<<<3'd2 )+$signed( -{ 2'b0,x368 }<<<3'd1 )+$signed( -{ 3'b0,x369 }<<<3'd2)+$signed( { 3'b0,x370 }<<<3'd2 )+$signed( { 3'b0,x371 }<<<3'd2 )+$signed( -{ 3'b0,x372 }<<<3'd2)+$signed( { 1'b0,x373 }  )+$signed( -{ 3'b0,x374 }<<<3'd2)+$signed( { 2'b0,x375 } <<<3'd1 )+$signed( -{ 3'b0,x376 }<<<3'd2)+$signed( { 2'b0,x377 } <<<3'd1 )+$signed( -{ 1'b0,x378 } )+$signed( { 1'b0,x379 }  )+$signed( { 2'b0,x382 } <<<3'd1 )+$signed( { 2'b0,x384 } <<<3'd1 )+$signed( { 3'b0,x385 }<<<3'd2 )+$signed( { 3'b0,x386 }<<<3'd2 )+$signed( -{ 2'b0,x388 }<<<3'd1 )+$signed( { 1'b0,x389 }  )+$signed( { 1'b0,x391 }  )+$signed( { 3'b0,x392 }<<<3'd2 )+$signed( -{ 3'b0,x393 }<<<3'd2)+$signed( { 2'b0,x395 } <<<3'd1 )+$signed( -{ 3'b0,x396 }<<<3'd2)+$signed( { 3'b0,x397 }<<<3'd2 )+$signed( -{ 1'b0,x398 } )+$signed( -{ 1'b0,x399 } )+$signed( -{ 2'b0,x401 }<<<3'd1 )+$signed( { 2'b0,x403 } <<<3'd1 )+$signed( -{ 2'b0,x404 }<<<3'd1 )+$signed( -{ 1'b0,x405 } )+$signed( { 1'b0,x406 }  )+$signed( { 1'b0,x407 }  )+$signed( -{ 1'b0,x408 } )+$signed( -{ 4'b0, x409 }<<<3'd3 )+$signed( -{ 1'b0,x410 } )+$signed( -{ 2'b0,x411 }<<<3'd1 )+$signed( { 1'b0,x412 }  )+$signed( -{ 1'b0,x413 } )+$signed( { 1'b0,x414 }  )+$signed( -{ 3'b0,x415 }<<<3'd2)+$signed( { 2'b0,x416 } <<<3'd1 )+$signed( -{ 2'b0,x417 }<<<3'd1 )+$signed( { 2'b0,x418 } <<<3'd1 )+$signed( { 2'b0,x419 } <<<3'd1 )+$signed( { 3'b0,x421 }<<<3'd2 )+$signed( -{ 3'b0,x422 }<<<3'd2)+$signed( { 2'b0,x423 } <<<3'd1 )+$signed( -{ 3'b0,x424 }<<<3'd2)+$signed( { 1'b0,x425 }  )+$signed( -{ 3'b0,x426 }<<<3'd2)+$signed( -{ 1'b0,x427 } )+$signed( -{ 2'b0,x428 }<<<3'd1 )+$signed( { 1'b0,x431 }  )+$signed( -{ 1'b0,x432 } )+$signed( { 1'b0,x433 }  )+$signed( -{ 1'b0,x434 } )+$signed( { 3'b0,x437 }<<<3'd2 )+$signed( -{ 3'b0,x439 }<<<3'd2)+$signed( -{ 4'b0, x442 }<<<3'd3 )+$signed( { 1'b0,x443 }  )+$signed( { 2'b0,x444 } <<<3'd1 )+$signed( -{ 3'b0,x445 }<<<3'd2)+$signed( -{ 1'b0,x446 } )+$signed( -{ 3'b0,x447 }<<<3'd2)+$signed( -{ 4'b0, x448 }<<<3'd3 )+$signed( -{ 2'b0,x449 }<<<3'd1 )+$signed( -{ 4'b0, x450 }<<<3'd3 )+$signed( { 3'b0,x451 }<<<3'd2 )+$signed( { 2'b0,x452 } <<<3'd1 )+$signed( { 1'b0,x453 }  )+$signed( -{ 3'b0,x454 }<<<3'd2)+$signed( { 1'b0,x455 }  )+$signed( { 2'b0,x457 } <<<3'd1 )+$signed( -{ 3'b0,x458 }<<<3'd2)+$signed( -{ 3'b0,x459 }<<<3'd2)+$signed( -{ 4'b0, x461 }<<<3'd3 )+$signed( { 2'b0,x462 } <<<3'd1 )+$signed( -{ 4'b0, x463 }<<<3'd3 )+$signed( { 3'b0,x464 }<<<3'd2 )+$signed( { 2'b0,x465 } <<<3'd1 )+$signed( -{ 2'b0,x466 }<<<3'd1 )+$signed( -{ 4'b0, x467 }<<<3'd3 )+$signed( -{ 2'b0,x468 }<<<3'd1 )+$signed( { 2'b0,x469 } <<<3'd1 )+$signed( { 3'b0,x470 }<<<3'd2 )+$signed( { 3'b0,x471 }<<<3'd2 )+$signed( -{ 3'b0,x472 }<<<3'd2)+$signed( -{ 1'b0,x473 } )+$signed( -{ 3'b0,x474 }<<<3'd2)+$signed( { 2'b0,x475 } <<<3'd1 )+$signed( -{ 3'b0,x476 }<<<3'd2)+$signed( -{ 2'b0,x477 }<<<3'd1 )+$signed( { 2'b0,x478 } <<<3'd1 )+$signed( { 3'b0,x479 }<<<3'd2 )+$signed( -{ 2'b0,x480 }<<<3'd1 )+$signed( { 1'b0,x481 }  )+$signed( { 1'b0,x482 }  )+$signed( { 1'b0,x483 }  )+$signed( -{ 3'b0,x484 }<<<3'd2)+$signed( { 1'b0,x485 }  )+$signed( { 3'b0,x487 }<<<3'd2 )+$signed( { 1'b0,x489 }  )+$signed( -{ 2'b0,x490 }<<<3'd1 )+$signed( { 1'b0,x491 }  )+$signed( { 3'b0,x492 }<<<3'd2 )+$signed( { 1'b0,x493 }  )+$signed( { 3'b0,x494 }<<<3'd2 )+$signed( -{ 1'b0,x495 } )+$signed(13'd8);
assign y9=temp_y[9][13] ==1'b1 ? 6'd0 :  
    temp_y[9][10] ==1'b1 ? 6'd63 : 
    temp_y[9][3]==1'b1 ? temp_y[9][9:4]+1'b1 : temp_y[9][9:4];
assign temp_y[10] = 
+$signed( -{ 3'b0,x0 }<<<3'd2)+$signed( -{ 1'b0,x1 } )+$signed( { 2'b0,x2 } <<<3'd1 )+$signed( { 1'b0,x3 }  )+$signed( -{ 2'b0,x4 }<<<3'd1 )+$signed( -{ 1'b0,x5 } )+$signed( { 3'b0,x6 }<<<3'd2 )+$signed( { 3'b0,x7 }<<<3'd2 )+$signed( { 3'b0,x8 }<<<3'd2 )+$signed( -{ 2'b0,x9 }<<<3'd1 )+$signed( -{ 1'b0,x10 } )+$signed( -{ 2'b0,x12 }<<<3'd1 )+$signed( -{ 2'b0,x13 }<<<3'd1 )+$signed( { 2'b0,x14 } <<<3'd1 )+$signed( { 2'b0,x15 } <<<3'd1 )+$signed( { 2'b0,x17 } <<<3'd1 )+$signed( -{ 2'b0,x18 }<<<3'd1 )+$signed( -{ 2'b0,x19 }<<<3'd1 )+$signed( -{ 1'b0,x20 } )+$signed( { 2'b0,x21 } <<<3'd1 )+$signed( { 2'b0,x22 } <<<3'd1 )+$signed( -{ 2'b0,x23 }<<<3'd1 )+$signed( -{ 1'b0,x24 } )+$signed( { 1'b0,x25 }  )+$signed( { 3'b0,x26 }<<<3'd2 )+$signed( -{ 3'b0,x27 }<<<3'd2)+$signed( { 3'b0,x28 }<<<3'd2 )+$signed( { 1'b0,x29 }  )+$signed( { 3'b0,x30 }<<<3'd2 )+$signed( -{ 1'b0,x31 } )+$signed( { 2'b0,x32 } <<<3'd1 )+$signed( -{ 1'b0,x33 } )+$signed( -{ 1'b0,x34 } )+$signed( { 1'b0,x35 }  )+$signed( -{ 3'b0,x36 }<<<3'd2)+$signed( -{ 2'b0,x37 }<<<3'd1 )+$signed( -{ 2'b0,x38 }<<<3'd1 )+$signed( { 1'b0,x40 }  )+$signed( -{ 1'b0,x41 } )+$signed( { 3'b0,x43 }<<<3'd2 )+$signed( { 2'b0,x44 } <<<3'd1 )+$signed( -{ 3'b0,x45 }<<<3'd2)+$signed( { 2'b0,x48 } <<<3'd1 )+$signed( -{ 1'b0,x49 } )+$signed( { 3'b0,x50 }<<<3'd2 )+$signed( -{ 2'b0,x52 }<<<3'd1 )+$signed( { 2'b0,x54 } <<<3'd1 )+$signed( -{ 2'b0,x55 }<<<3'd1 )+$signed( { 2'b0,x56 } <<<3'd1 )+$signed( -{ 1'b0,x57 } )+$signed( { 3'b0,x58 }<<<3'd2 )+$signed( { 1'b0,x59 }  )+$signed( { 1'b0,x60 }  )+$signed( -{ 1'b0,x61 } )+$signed( { 2'b0,x62 } <<<3'd1 )+$signed( { 2'b0,x63 } <<<3'd1 )+$signed( -{ 2'b0,x64 }<<<3'd1 )+$signed( { 2'b0,x65 } <<<3'd1 )+$signed( -{ 2'b0,x66 }<<<3'd1 )+$signed( -{ 1'b0,x67 } )+$signed( { 2'b0,x68 } <<<3'd1 )+$signed( { 3'b0,x69 }<<<3'd2 )+$signed( -{ 1'b0,x70 } )+$signed( { 2'b0,x71 } <<<3'd1 )+$signed( -{ 2'b0,x72 }<<<3'd1 )+$signed( { 1'b0,x73 }  )+$signed( { 3'b0,x75 }<<<3'd2 )+$signed( { 3'b0,x76 }<<<3'd2 )+$signed( { 2'b0,x77 } <<<3'd1 )+$signed( { 3'b0,x78 }<<<3'd2 )+$signed( -{ 2'b0,x80 }<<<3'd1 )+$signed( -{ 1'b0,x81 } )+$signed( -{ 1'b0,x82 } )+$signed( { 3'b0,x83 }<<<3'd2 )+$signed( -{ 3'b0,x84 }<<<3'd2)+$signed( -{ 3'b0,x85 }<<<3'd2)+$signed( -{ 2'b0,x86 }<<<3'd1 )+$signed( -{ 2'b0,x87 }<<<3'd1 )+$signed( -{ 1'b0,x88 } )+$signed( { 3'b0,x89 }<<<3'd2 )+$signed( { 3'b0,x90 }<<<3'd2 )+$signed( -{ 3'b0,x91 }<<<3'd2)+$signed( { 1'b0,x92 }  )+$signed( { 2'b0,x93 } <<<3'd1 )+$signed( { 3'b0,x94 }<<<3'd2 )+$signed( { 1'b0,x95 }  )+$signed( { 2'b0,x96 } <<<3'd1 )+$signed( { 1'b0,x97 }  )+$signed( { 3'b0,x98 }<<<3'd2 )+$signed( -{ 4'b0, x99 }<<<3'd3 )+$signed( -{ 3'b0,x100 }<<<3'd2)+$signed( -{ 3'b0,x101 }<<<3'd2)+$signed( -{ 3'b0,x102 }<<<3'd2)+$signed( -{ 2'b0,x103 }<<<3'd1 )+$signed( { 3'b0,x104 }<<<3'd2 )+$signed( -{ 2'b0,x105 }<<<3'd1 )+$signed( { 1'b0,x106 }  )+$signed( -{ 1'b0,x107 } )+$signed( -{ 1'b0,x108 } )+$signed( -{ 3'b0,x109 }<<<3'd2)+$signed( { 1'b0,x110 }  )+$signed( { 2'b0,x111 } <<<3'd1 )+$signed( { 4'b0,x112 }<<<3'd3 )+$signed( { 2'b0,x114 } <<<3'd1 )+$signed( { 4'b0,x116 }<<<3'd3 )+$signed( -{ 3'b0,x117 }<<<3'd2)+$signed( -{ 3'b0,x118 }<<<3'd2)+$signed( -{ 3'b0,x119 }<<<3'd2)+$signed( -{ 3'b0,x120 }<<<3'd2)+$signed( -{ 1'b0,x121 } )+$signed( -{ 2'b0,x122 }<<<3'd1 )+$signed( { 1'b0,x123 }  )+$signed( -{ 2'b0,x124 }<<<3'd1 )+$signed( -{ 2'b0,x125 }<<<3'd1 )+$signed( -{ 2'b0,x126 }<<<3'd1 )+$signed( { 2'b0,x127 } <<<3'd1 )+$signed( { 2'b0,x128 } <<<3'd1 )+$signed( { 4'b0,x129 }<<<3'd3 )+$signed( { 2'b0,x130 } <<<3'd1 )+$signed( -{ 2'b0,x131 }<<<3'd1 )+$signed( -{ 2'b0,x133 }<<<3'd1 )+$signed( { 1'b0,x134 }  )+$signed( -{ 2'b0,x135 }<<<3'd1 )+$signed( { 1'b0,x136 }  )+$signed( { 1'b0,x137 }  )+$signed( -{ 3'b0,x138 }<<<3'd2)+$signed( -{ 2'b0,x139 }<<<3'd1 )+$signed( -{ 3'b0,x140 }<<<3'd2)+$signed( { 2'b0,x141 } <<<3'd1 )+$signed( { 2'b0,x142 } <<<3'd1 )+$signed( { 3'b0,x143 }<<<3'd2 )+$signed( -{ 3'b0,x144 }<<<3'd2)+$signed( { 2'b0,x145 } <<<3'd1 )+$signed( -{ 3'b0,x146 }<<<3'd2)+$signed( -{ 1'b0,x147 } )+$signed( -{ 1'b0,x148 } )+$signed( -{ 2'b0,x150 }<<<3'd1 )+$signed( { 2'b0,x151 } <<<3'd1 )+$signed( { 1'b0,x152 }  )+$signed( { 2'b0,x154 } <<<3'd1 )+$signed( -{ 2'b0,x156 }<<<3'd1 )+$signed( -{ 3'b0,x157 }<<<3'd2)+$signed( { 1'b0,x158 }  )+$signed( -{ 2'b0,x159 }<<<3'd1 )+$signed( -{ 1'b0,x160 } )+$signed( { 3'b0,x161 }<<<3'd2 )+$signed( -{ 3'b0,x162 }<<<3'd2)+$signed( { 2'b0,x163 } <<<3'd1 )+$signed( -{ 1'b0,x164 } )+$signed( { 2'b0,x165 } <<<3'd1 )+$signed( { 2'b0,x166 } <<<3'd1 )+$signed( { 3'b0,x168 }<<<3'd2 )+$signed( -{ 1'b0,x169 } )+$signed( { 3'b0,x170 }<<<3'd2 )+$signed( -{ 3'b0,x171 }<<<3'd2)+$signed( -{ 3'b0,x175 }<<<3'd2)+$signed( { 3'b0,x176 }<<<3'd2 )+$signed( -{ 3'b0,x177 }<<<3'd2)+$signed( -{ 1'b0,x178 } )+$signed( -{ 2'b0,x179 }<<<3'd1 )+$signed( { 1'b0,x180 }  )+$signed( { 1'b0,x181 }  )+$signed( -{ 2'b0,x182 }<<<3'd1 )+$signed( -{ 3'b0,x183 }<<<3'd2)+$signed( { 3'b0,x184 }<<<3'd2 )+$signed( { 3'b0,x186 }<<<3'd2 )+$signed( -{ 1'b0,x187 } )+$signed( { 3'b0,x188 }<<<3'd2 )+$signed( -{ 4'b0, x189 }<<<3'd3 )+$signed( { 1'b0,x190 }  )+$signed( { 1'b0,x191 }  )+$signed( -{ 2'b0,x192 }<<<3'd1 )+$signed( -{ 3'b0,x193 }<<<3'd2)+$signed( -{ 1'b0,x194 } )+$signed( -{ 3'b0,x195 }<<<3'd2)+$signed( { 3'b0,x196 }<<<3'd2 )+$signed( { 1'b0,x197 }  )+$signed( { 1'b0,x201 }  )+$signed( -{ 1'b0,x202 } )+$signed( { 3'b0,x203 }<<<3'd2 )+$signed( -{ 2'b0,x205 }<<<3'd1 )+$signed( { 3'b0,x206 }<<<3'd2 )+$signed( -{ 2'b0,x207 }<<<3'd1 )+$signed( { 1'b0,x208 }  )+$signed( { 2'b0,x209 } <<<3'd1 )+$signed( -{ 2'b0,x210 }<<<3'd1 )+$signed( -{ 3'b0,x211 }<<<3'd2)+$signed( { 3'b0,x212 }<<<3'd2 )+$signed( { 1'b0,x213 }  )+$signed( -{ 2'b0,x214 }<<<3'd1 )+$signed( { 3'b0,x215 }<<<3'd2 )+$signed( { 3'b0,x216 }<<<3'd2 )+$signed( { 3'b0,x217 }<<<3'd2 )+$signed( -{ 2'b0,x218 }<<<3'd1 )+$signed( -{ 3'b0,x219 }<<<3'd2)+$signed( { 2'b0,x220 } <<<3'd1 )+$signed( -{ 2'b0,x221 }<<<3'd1 )+$signed( { 2'b0,x223 } <<<3'd1 )+$signed( { 2'b0,x224 } <<<3'd1 )+$signed( -{ 1'b0,x225 } )+$signed( -{ 3'b0,x226 }<<<3'd2)+$signed( { 2'b0,x227 } <<<3'd1 )+$signed( { 1'b0,x228 }  )+$signed( { 2'b0,x229 } <<<3'd1 )+$signed( { 3'b0,x231 }<<<3'd2 )+$signed( { 2'b0,x232 } <<<3'd1 )+$signed( { 3'b0,x233 }<<<3'd2 )+$signed( { 1'b0,x234 }  )+$signed( { 3'b0,x235 }<<<3'd2 )+$signed( -{ 2'b0,x236 }<<<3'd1 )+$signed( -{ 2'b0,x237 }<<<3'd1 )+$signed( { 3'b0,x238 }<<<3'd2 )+$signed( -{ 1'b0,x239 } )+$signed( { 3'b0,x240 }<<<3'd2 )+$signed( { 2'b0,x241 } <<<3'd1 )+$signed( -{ 3'b0,x243 }<<<3'd2)+$signed( -{ 2'b0,x244 }<<<3'd1 )+$signed( { 1'b0,x245 }  )+$signed( -{ 2'b0,x246 }<<<3'd1 )+$signed( { 1'b0,x247 }  )+$signed( -{ 1'b0,x248 } )+$signed( -{ 2'b0,x249 }<<<3'd1 )+$signed( { 3'b0,x250 }<<<3'd2 )+$signed( { 3'b0,x251 }<<<3'd2 )+$signed( -{ 2'b0,x252 }<<<3'd1 )+$signed( { 3'b0,x253 }<<<3'd2 )+$signed( -{ 3'b0,x255 }<<<3'd2)+$signed( { 2'b0,x256 } <<<3'd1 )+$signed( -{ 1'b0,x257 } )+$signed( { 3'b0,x258 }<<<3'd2 )+$signed( { 2'b0,x259 } <<<3'd1 )+$signed( { 2'b0,x260 } <<<3'd1 )+$signed( -{ 3'b0,x261 }<<<3'd2)+$signed( -{ 3'b0,x262 }<<<3'd2)+$signed( -{ 3'b0,x264 }<<<3'd2)+$signed( -{ 1'b0,x266 } )+$signed( -{ 1'b0,x267 } )+$signed( -{ 1'b0,x268 } )+$signed( { 2'b0,x269 } <<<3'd1 )+$signed( { 3'b0,x270 }<<<3'd2 )+$signed( { 3'b0,x271 }<<<3'd2 )+$signed( -{ 2'b0,x273 }<<<3'd1 )+$signed( { 1'b0,x274 }  )+$signed( -{ 3'b0,x275 }<<<3'd2)+$signed( { 1'b0,x276 }  )+$signed( { 1'b0,x277 }  )+$signed( { 2'b0,x278 } <<<3'd1 )+$signed( -{ 2'b0,x279 }<<<3'd1 )+$signed( -{ 3'b0,x280 }<<<3'd2)+$signed( { 1'b0,x281 }  )+$signed( { 2'b0,x282 } <<<3'd1 )+$signed( -{ 2'b0,x283 }<<<3'd1 )+$signed( -{ 1'b0,x284 } )+$signed( -{ 2'b0,x285 }<<<3'd1 )+$signed( { 2'b0,x286 } <<<3'd1 )+$signed( { 2'b0,x287 } <<<3'd1 )+$signed( -{ 2'b0,x288 }<<<3'd1 )+$signed( { 2'b0,x290 } <<<3'd1 )+$signed( -{ 2'b0,x291 }<<<3'd1 )+$signed( { 3'b0,x292 }<<<3'd2 )+$signed( -{ 3'b0,x293 }<<<3'd2)+$signed( { 2'b0,x294 } <<<3'd1 )+$signed( { 2'b0,x295 } <<<3'd1 )+$signed( { 3'b0,x296 }<<<3'd2 )+$signed( { 2'b0,x297 } <<<3'd1 )+$signed( -{ 1'b0,x298 } )+$signed( { 2'b0,x299 } <<<3'd1 )+$signed( -{ 2'b0,x300 }<<<3'd1 )+$signed( -{ 3'b0,x301 }<<<3'd2)+$signed( { 3'b0,x303 }<<<3'd2 )+$signed( { 2'b0,x304 } <<<3'd1 )+$signed( { 2'b0,x305 } <<<3'd1 )+$signed( { 1'b0,x306 }  )+$signed( -{ 2'b0,x307 }<<<3'd1 )+$signed( -{ 2'b0,x308 }<<<3'd1 )+$signed( { 2'b0,x309 } <<<3'd1 )+$signed( -{ 1'b0,x310 } )+$signed( -{ 2'b0,x311 }<<<3'd1 )+$signed( -{ 1'b0,x312 } )+$signed( -{ 1'b0,x313 } )+$signed( { 2'b0,x314 } <<<3'd1 )+$signed( { 3'b0,x316 }<<<3'd2 )+$signed( -{ 3'b0,x317 }<<<3'd2)+$signed( -{ 2'b0,x318 }<<<3'd1 )+$signed( -{ 2'b0,x319 }<<<3'd1 )+$signed( { 1'b0,x321 }  )+$signed( { 2'b0,x322 } <<<3'd1 )+$signed( -{ 3'b0,x323 }<<<3'd2)+$signed( -{ 1'b0,x324 } )+$signed( -{ 1'b0,x325 } )+$signed( { 3'b0,x326 }<<<3'd2 )+$signed( -{ 2'b0,x328 }<<<3'd1 )+$signed( { 2'b0,x329 } <<<3'd1 )+$signed( -{ 2'b0,x330 }<<<3'd1 )+$signed( -{ 3'b0,x331 }<<<3'd2)+$signed( -{ 2'b0,x332 }<<<3'd1 )+$signed( { 2'b0,x333 } <<<3'd1 )+$signed( { 2'b0,x334 } <<<3'd1 )+$signed( { 2'b0,x337 } <<<3'd1 )+$signed( { 1'b0,x338 }  )+$signed( -{ 1'b0,x341 } )+$signed( { 4'b0,x342 }<<<3'd3 )+$signed( -{ 2'b0,x343 }<<<3'd1 )+$signed( { 2'b0,x344 } <<<3'd1 )+$signed( -{ 2'b0,x345 }<<<3'd1 )+$signed( { 2'b0,x346 } <<<3'd1 )+$signed( -{ 1'b0,x347 } )+$signed( { 3'b0,x348 }<<<3'd2 )+$signed( { 1'b0,x349 }  )+$signed( { 1'b0,x350 }  )+$signed( { 3'b0,x351 }<<<3'd2 )+$signed( { 1'b0,x352 }  )+$signed( { 1'b0,x353 }  )+$signed( { 1'b0,x354 }  )+$signed( { 3'b0,x355 }<<<3'd2 )+$signed( -{ 2'b0,x356 }<<<3'd1 )+$signed( -{ 3'b0,x358 }<<<3'd2)+$signed( { 1'b0,x359 }  )+$signed( -{ 1'b0,x360 } )+$signed( { 1'b0,x361 }  )+$signed( { 3'b0,x362 }<<<3'd2 )+$signed( -{ 2'b0,x363 }<<<3'd1 )+$signed( -{ 1'b0,x364 } )+$signed( { 3'b0,x365 }<<<3'd2 )+$signed( -{ 2'b0,x367 }<<<3'd1 )+$signed( -{ 1'b0,x368 } )+$signed( -{ 3'b0,x369 }<<<3'd2)+$signed( { 2'b0,x370 } <<<3'd1 )+$signed( -{ 3'b0,x371 }<<<3'd2)+$signed( { 2'b0,x374 } <<<3'd1 )+$signed( { 3'b0,x375 }<<<3'd2 )+$signed( { 3'b0,x377 }<<<3'd2 )+$signed( { 2'b0,x378 } <<<3'd1 )+$signed( { 1'b0,x379 }  )+$signed( -{ 1'b0,x380 } )+$signed( { 4'b0,x381 }<<<3'd3 )+$signed( -{ 3'b0,x382 }<<<3'd2)+$signed( -{ 3'b0,x383 }<<<3'd2)+$signed( -{ 3'b0,x384 }<<<3'd2)+$signed( { 2'b0,x385 } <<<3'd1 )+$signed( -{ 1'b0,x386 } )+$signed( -{ 1'b0,x387 } )+$signed( -{ 2'b0,x388 }<<<3'd1 )+$signed( { 2'b0,x389 } <<<3'd1 )+$signed( { 3'b0,x390 }<<<3'd2 )+$signed( { 3'b0,x391 }<<<3'd2 )+$signed( -{ 2'b0,x392 }<<<3'd1 )+$signed( -{ 1'b0,x393 } )+$signed( { 2'b0,x394 } <<<3'd1 )+$signed( -{ 2'b0,x395 }<<<3'd1 )+$signed( { 1'b0,x396 }  )+$signed( { 2'b0,x397 } <<<3'd1 )+$signed( -{ 2'b0,x398 }<<<3'd1 )+$signed( { 1'b0,x399 }  )+$signed( { 1'b0,x401 }  )+$signed( { 2'b0,x402 } <<<3'd1 )+$signed( { 2'b0,x404 } <<<3'd1 )+$signed( { 2'b0,x405 } <<<3'd1 )+$signed( -{ 2'b0,x406 }<<<3'd1 )+$signed( { 3'b0,x407 }<<<3'd2 )+$signed( -{ 1'b0,x408 } )+$signed( { 3'b0,x409 }<<<3'd2 )+$signed( -{ 2'b0,x410 }<<<3'd1 )+$signed( -{ 2'b0,x411 }<<<3'd1 )+$signed( -{ 2'b0,x415 }<<<3'd1 )+$signed( -{ 4'b0, x416 }<<<3'd3 )+$signed( { 3'b0,x417 }<<<3'd2 )+$signed( { 1'b0,x420 }  )+$signed( -{ 2'b0,x421 }<<<3'd1 )+$signed( -{ 2'b0,x422 }<<<3'd1 )+$signed( { 2'b0,x423 } <<<3'd1 )+$signed( -{ 1'b0,x424 } )+$signed( { 2'b0,x425 } <<<3'd1 )+$signed( -{ 2'b0,x426 }<<<3'd1 )+$signed( { 2'b0,x427 } <<<3'd1 )+$signed( -{ 2'b0,x428 }<<<3'd1 )+$signed( -{ 1'b0,x429 } )+$signed( { 3'b0,x430 }<<<3'd2 )+$signed( { 2'b0,x431 } <<<3'd1 )+$signed( -{ 3'b0,x432 }<<<3'd2)+$signed( -{ 1'b0,x433 } )+$signed( -{ 3'b0,x434 }<<<3'd2)+$signed( -{ 3'b0,x435 }<<<3'd2)+$signed( -{ 2'b0,x436 }<<<3'd1 )+$signed( -{ 1'b0,x437 } )+$signed( -{ 1'b0,x439 } )+$signed( { 2'b0,x440 } <<<3'd1 )+$signed( -{ 2'b0,x441 }<<<3'd1 )+$signed( -{ 2'b0,x442 }<<<3'd1 )+$signed( { 3'b0,x443 }<<<3'd2 )+$signed( { 3'b0,x445 }<<<3'd2 )+$signed( -{ 2'b0,x446 }<<<3'd1 )+$signed( { 1'b0,x447 }  )+$signed( { 3'b0,x448 }<<<3'd2 )+$signed( -{ 2'b0,x449 }<<<3'd1 )+$signed( { 2'b0,x451 } <<<3'd1 )+$signed( -{ 2'b0,x452 }<<<3'd1 )+$signed( -{ 1'b0,x454 } )+$signed( -{ 2'b0,x455 }<<<3'd1 )+$signed( -{ 2'b0,x456 }<<<3'd1 )+$signed( -{ 1'b0,x457 } )+$signed( { 1'b0,x459 }  )+$signed( -{ 2'b0,x460 }<<<3'd1 )+$signed( { 2'b0,x461 } <<<3'd1 )+$signed( { 1'b0,x462 }  )+$signed( -{ 1'b0,x463 } )+$signed( -{ 2'b0,x466 }<<<3'd1 )+$signed( -{ 3'b0,x468 }<<<3'd2)+$signed( { 1'b0,x471 }  )+$signed( -{ 3'b0,x472 }<<<3'd2)+$signed( { 1'b0,x474 }  )+$signed( { 2'b0,x475 } <<<3'd1 )+$signed( { 1'b0,x476 }  )+$signed( { 3'b0,x478 }<<<3'd2 )+$signed( { 1'b0,x480 }  )+$signed( { 3'b0,x481 }<<<3'd2 )+$signed( { 1'b0,x482 }  )+$signed( -{ 1'b0,x483 } )+$signed( { 3'b0,x484 }<<<3'd2 )+$signed( -{ 2'b0,x485 }<<<3'd1 )+$signed( -{ 2'b0,x486 }<<<3'd1 )+$signed( { 2'b0,x487 } <<<3'd1 )+$signed( { 1'b0,x488 }  )+$signed( { 1'b0,x489 }  )+$signed( { 2'b0,x490 } <<<3'd1 )+$signed( -{ 2'b0,x491 }<<<3'd1 )+$signed( { 2'b0,x492 } <<<3'd1 )+$signed( -{ 2'b0,x493 }<<<3'd1 )+$signed( { 1'b0,x494 }  )+$signed( -{ 1'b0,x495 } )+$signed(13'd56);
assign y10=temp_y[10][13] ==1'b1 ? 6'd0 :  
    temp_y[10][10] ==1'b1 ? 6'd63 : 
    temp_y[10][3]==1'b1 ? temp_y[10][9:4]+1'b1 : temp_y[10][9:4];
assign temp_y[11] = 
+$signed( -{ 3'b0,x0 }<<<3'd2)+$signed( { 2'b0,x2 } <<<3'd1 )+$signed( { 1'b0,x3 }  )+$signed( -{ 1'b0,x4 } )+$signed( { 2'b0,x6 } <<<3'd1 )+$signed( -{ 1'b0,x7 } )+$signed( { 1'b0,x8 }  )+$signed( { 2'b0,x9 } <<<3'd1 )+$signed( -{ 3'b0,x10 }<<<3'd2)+$signed( -{ 1'b0,x11 } )+$signed( -{ 3'b0,x12 }<<<3'd2)+$signed( -{ 1'b0,x13 } )+$signed( -{ 1'b0,x14 } )+$signed( { 2'b0,x15 } <<<3'd1 )+$signed( { 2'b0,x16 } <<<3'd1 )+$signed( { 3'b0,x18 }<<<3'd2 )+$signed( -{ 2'b0,x20 }<<<3'd1 )+$signed( -{ 1'b0,x21 } )+$signed( { 3'b0,x22 }<<<3'd2 )+$signed( -{ 1'b0,x23 } )+$signed( -{ 1'b0,x24 } )+$signed( -{ 1'b0,x25 } )+$signed( -{ 2'b0,x26 }<<<3'd1 )+$signed( { 1'b0,x27 }  )+$signed( { 3'b0,x30 }<<<3'd2 )+$signed( -{ 3'b0,x32 }<<<3'd2)+$signed( -{ 2'b0,x33 }<<<3'd1 )+$signed( { 1'b0,x34 }  )+$signed( -{ 1'b0,x35 } )+$signed( { 1'b0,x36 }  )+$signed( { 2'b0,x37 } <<<3'd1 )+$signed( -{ 1'b0,x38 } )+$signed( -{ 2'b0,x39 }<<<3'd1 )+$signed( { 2'b0,x40 } <<<3'd1 )+$signed( -{ 1'b0,x43 } )+$signed( -{ 2'b0,x44 }<<<3'd1 )+$signed( -{ 2'b0,x46 }<<<3'd1 )+$signed( { 2'b0,x47 } <<<3'd1 )+$signed( { 3'b0,x48 }<<<3'd2 )+$signed( -{ 1'b0,x49 } )+$signed( { 1'b0,x50 }  )+$signed( { 2'b0,x51 } <<<3'd1 )+$signed( { 3'b0,x52 }<<<3'd2 )+$signed( -{ 1'b0,x53 } )+$signed( { 1'b0,x54 }  )+$signed( { 2'b0,x55 } <<<3'd1 )+$signed( { 2'b0,x56 } <<<3'd1 )+$signed( -{ 1'b0,x57 } )+$signed( { 1'b0,x58 }  )+$signed( -{ 1'b0,x59 } )+$signed( -{ 2'b0,x61 }<<<3'd1 )+$signed( { 1'b0,x62 }  )+$signed( -{ 2'b0,x63 }<<<3'd1 )+$signed( -{ 3'b0,x64 }<<<3'd2)+$signed( -{ 1'b0,x65 } )+$signed( { 1'b0,x67 }  )+$signed( { 1'b0,x68 }  )+$signed( -{ 2'b0,x69 }<<<3'd1 )+$signed( { 2'b0,x70 } <<<3'd1 )+$signed( -{ 2'b0,x73 }<<<3'd1 )+$signed( -{ 1'b0,x74 } )+$signed( -{ 1'b0,x75 } )+$signed( { 1'b0,x76 }  )+$signed( -{ 1'b0,x77 } )+$signed( { 3'b0,x78 }<<<3'd2 )+$signed( -{ 2'b0,x79 }<<<3'd1 )+$signed( { 2'b0,x80 } <<<3'd1 )+$signed( { 1'b0,x81 }  )+$signed( -{ 3'b0,x82 }<<<3'd2)+$signed( { 1'b0,x85 }  )+$signed( { 1'b0,x86 }  )+$signed( { 1'b0,x87 }  )+$signed( { 1'b0,x88 }  )+$signed( -{ 1'b0,x89 } )+$signed( { 3'b0,x90 }<<<3'd2 )+$signed( { 3'b0,x91 }<<<3'd2 )+$signed( -{ 2'b0,x92 }<<<3'd1 )+$signed( -{ 2'b0,x93 }<<<3'd1 )+$signed( { 4'b0,x94 }<<<3'd3 )+$signed( -{ 3'b0,x95 }<<<3'd2)+$signed( -{ 4'b0, x96 }<<<3'd3 )+$signed( { 2'b0,x97 } <<<3'd1 )+$signed( -{ 3'b0,x98 }<<<3'd2)+$signed( { 2'b0,x99 } <<<3'd1 )+$signed( { 3'b0,x100 }<<<3'd2 )+$signed( { 3'b0,x101 }<<<3'd2 )+$signed( { 3'b0,x102 }<<<3'd2 )+$signed( { 2'b0,x103 } <<<3'd1 )+$signed( -{ 3'b0,x104 }<<<3'd2)+$signed( { 2'b0,x105 } <<<3'd1 )+$signed( { 2'b0,x106 } <<<3'd1 )+$signed( { 1'b0,x107 }  )+$signed( { 3'b0,x108 }<<<3'd2 )+$signed( { 3'b0,x109 }<<<3'd2 )+$signed( -{ 2'b0,x110 }<<<3'd1 )+$signed( -{ 3'b0,x111 }<<<3'd2)+$signed( { 3'b0,x112 }<<<3'd2 )+$signed( -{ 1'b0,x113 } )+$signed( -{ 4'b0, x114 }<<<3'd3 )+$signed( { 3'b0,x115 }<<<3'd2 )+$signed( -{ 3'b0,x116 }<<<3'd2)+$signed( -{ 2'b0,x117 }<<<3'd1 )+$signed( { 3'b0,x118 }<<<3'd2 )+$signed( { 3'b0,x119 }<<<3'd2 )+$signed( { 3'b0,x120 }<<<3'd2 )+$signed( { 3'b0,x121 }<<<3'd2 )+$signed( -{ 1'b0,x122 } )+$signed( { 1'b0,x123 }  )+$signed( { 2'b0,x124 } <<<3'd1 )+$signed( { 2'b0,x125 } <<<3'd1 )+$signed( -{ 2'b0,x126 }<<<3'd1 )+$signed( { 1'b0,x127 }  )+$signed( { 1'b0,x128 }  )+$signed( -{ 2'b0,x129 }<<<3'd1 )+$signed( { 1'b0,x130 }  )+$signed( { 3'b0,x131 }<<<3'd2 )+$signed( -{ 2'b0,x132 }<<<3'd1 )+$signed( { 1'b0,x133 }  )+$signed( -{ 1'b0,x134 } )+$signed( { 3'b0,x135 }<<<3'd2 )+$signed( -{ 3'b0,x136 }<<<3'd2)+$signed( { 3'b0,x138 }<<<3'd2 )+$signed( { 2'b0,x139 } <<<3'd1 )+$signed( -{ 1'b0,x140 } )+$signed( { 1'b0,x141 }  )+$signed( { 2'b0,x142 } <<<3'd1 )+$signed( -{ 2'b0,x143 }<<<3'd1 )+$signed( -{ 1'b0,x144 } )+$signed( -{ 2'b0,x145 }<<<3'd1 )+$signed( -{ 1'b0,x146 } )+$signed( { 3'b0,x147 }<<<3'd2 )+$signed( { 2'b0,x148 } <<<3'd1 )+$signed( { 2'b0,x149 } <<<3'd1 )+$signed( { 2'b0,x150 } <<<3'd1 )+$signed( { 3'b0,x152 }<<<3'd2 )+$signed( -{ 1'b0,x153 } )+$signed( -{ 3'b0,x154 }<<<3'd2)+$signed( { 2'b0,x155 } <<<3'd1 )+$signed( { 2'b0,x156 } <<<3'd1 )+$signed( -{ 1'b0,x157 } )+$signed( { 2'b0,x158 } <<<3'd1 )+$signed( -{ 1'b0,x159 } )+$signed( { 1'b0,x160 }  )+$signed( -{ 1'b0,x161 } )+$signed( { 1'b0,x162 }  )+$signed( { 4'b0,x163 }<<<3'd3 )+$signed( { 3'b0,x164 }<<<3'd2 )+$signed( { 1'b0,x165 }  )+$signed( { 1'b0,x166 }  )+$signed( -{ 2'b0,x167 }<<<3'd1 )+$signed( -{ 3'b0,x168 }<<<3'd2)+$signed( { 3'b0,x169 }<<<3'd2 )+$signed( { 1'b0,x170 }  )+$signed( { 3'b0,x171 }<<<3'd2 )+$signed( { 3'b0,x172 }<<<3'd2 )+$signed( { 1'b0,x173 }  )+$signed( { 2'b0,x174 } <<<3'd1 )+$signed( { 3'b0,x175 }<<<3'd2 )+$signed( { 2'b0,x176 } <<<3'd1 )+$signed( -{ 1'b0,x177 } )+$signed( { 3'b0,x178 }<<<3'd2 )+$signed( -{ 2'b0,x179 }<<<3'd1 )+$signed( { 2'b0,x180 } <<<3'd1 )+$signed( { 4'b0,x181 }<<<3'd3 )+$signed( { 1'b0,x183 }  )+$signed( { 2'b0,x184 } <<<3'd1 )+$signed( -{ 2'b0,x185 }<<<3'd1 )+$signed( -{ 4'b0, x186 }<<<3'd3 )+$signed( { 1'b0,x188 }  )+$signed( { 3'b0,x189 }<<<3'd2 )+$signed( { 3'b0,x190 }<<<3'd2 )+$signed( { 3'b0,x191 }<<<3'd2 )+$signed( { 3'b0,x192 }<<<3'd2 )+$signed( { 3'b0,x193 }<<<3'd2 )+$signed( { 2'b0,x194 } <<<3'd1 )+$signed( { 2'b0,x195 } <<<3'd1 )+$signed( { 3'b0,x196 }<<<3'd2 )+$signed( -{ 3'b0,x197 }<<<3'd2)+$signed( { 2'b0,x199 } <<<3'd1 )+$signed( -{ 1'b0,x201 } )+$signed( -{ 2'b0,x202 }<<<3'd1 )+$signed( { 3'b0,x203 }<<<3'd2 )+$signed( { 1'b0,x204 }  )+$signed( { 2'b0,x205 } <<<3'd1 )+$signed( { 3'b0,x207 }<<<3'd2 )+$signed( -{ 2'b0,x208 }<<<3'd1 )+$signed( { 2'b0,x209 } <<<3'd1 )+$signed( { 3'b0,x210 }<<<3'd2 )+$signed( -{ 1'b0,x212 } )+$signed( { 1'b0,x213 }  )+$signed( { 1'b0,x214 }  )+$signed( -{ 2'b0,x215 }<<<3'd1 )+$signed( -{ 3'b0,x217 }<<<3'd2)+$signed( { 2'b0,x218 } <<<3'd1 )+$signed( -{ 3'b0,x220 }<<<3'd2)+$signed( { 1'b0,x221 }  )+$signed( { 3'b0,x222 }<<<3'd2 )+$signed( { 2'b0,x223 } <<<3'd1 )+$signed( { 3'b0,x224 }<<<3'd2 )+$signed( -{ 3'b0,x225 }<<<3'd2)+$signed( -{ 3'b0,x226 }<<<3'd2)+$signed( { 2'b0,x227 } <<<3'd1 )+$signed( -{ 1'b0,x228 } )+$signed( { 3'b0,x229 }<<<3'd2 )+$signed( { 2'b0,x230 } <<<3'd1 )+$signed( -{ 3'b0,x231 }<<<3'd2)+$signed( { 1'b0,x232 }  )+$signed( { 2'b0,x233 } <<<3'd1 )+$signed( -{ 3'b0,x234 }<<<3'd2)+$signed( -{ 1'b0,x235 } )+$signed( { 3'b0,x236 }<<<3'd2 )+$signed( { 1'b0,x238 }  )+$signed( -{ 2'b0,x239 }<<<3'd1 )+$signed( { 2'b0,x241 } <<<3'd1 )+$signed( { 2'b0,x242 } <<<3'd1 )+$signed( -{ 1'b0,x243 } )+$signed( -{ 3'b0,x244 }<<<3'd2)+$signed( { 2'b0,x245 } <<<3'd1 )+$signed( -{ 2'b0,x246 }<<<3'd1 )+$signed( -{ 2'b0,x247 }<<<3'd1 )+$signed( { 1'b0,x248 }  )+$signed( { 2'b0,x249 } <<<3'd1 )+$signed( -{ 2'b0,x251 }<<<3'd1 )+$signed( -{ 3'b0,x252 }<<<3'd2)+$signed( { 1'b0,x253 }  )+$signed( { 3'b0,x254 }<<<3'd2 )+$signed( { 2'b0,x255 } <<<3'd1 )+$signed( { 1'b0,x256 }  )+$signed( -{ 3'b0,x257 }<<<3'd2)+$signed( { 1'b0,x258 }  )+$signed( { 1'b0,x259 }  )+$signed( { 1'b0,x260 }  )+$signed( { 2'b0,x261 } <<<3'd1 )+$signed( { 1'b0,x263 }  )+$signed( { 2'b0,x266 } <<<3'd1 )+$signed( { 3'b0,x267 }<<<3'd2 )+$signed( { 1'b0,x268 }  )+$signed( -{ 2'b0,x269 }<<<3'd1 )+$signed( -{ 3'b0,x270 }<<<3'd2)+$signed( -{ 2'b0,x271 }<<<3'd1 )+$signed( -{ 1'b0,x272 } )+$signed( { 2'b0,x273 } <<<3'd1 )+$signed( -{ 3'b0,x274 }<<<3'd2)+$signed( { 3'b0,x275 }<<<3'd2 )+$signed( { 3'b0,x276 }<<<3'd2 )+$signed( { 1'b0,x277 }  )+$signed( { 3'b0,x278 }<<<3'd2 )+$signed( -{ 2'b0,x279 }<<<3'd1 )+$signed( -{ 3'b0,x280 }<<<3'd2)+$signed( { 2'b0,x281 } <<<3'd1 )+$signed( { 1'b0,x282 }  )+$signed( { 1'b0,x283 }  )+$signed( { 2'b0,x284 } <<<3'd1 )+$signed( { 2'b0,x286 } <<<3'd1 )+$signed( -{ 2'b0,x287 }<<<3'd1 )+$signed( -{ 1'b0,x288 } )+$signed( { 1'b0,x289 }  )+$signed( { 2'b0,x290 } <<<3'd1 )+$signed( -{ 2'b0,x291 }<<<3'd1 )+$signed( { 3'b0,x292 }<<<3'd2 )+$signed( -{ 1'b0,x293 } )+$signed( { 2'b0,x294 } <<<3'd1 )+$signed( { 3'b0,x295 }<<<3'd2 )+$signed( -{ 1'b0,x296 } )+$signed( -{ 1'b0,x297 } )+$signed( { 1'b0,x298 }  )+$signed( -{ 2'b0,x299 }<<<3'd1 )+$signed( -{ 2'b0,x300 }<<<3'd1 )+$signed( { 2'b0,x301 } <<<3'd1 )+$signed( { 2'b0,x302 } <<<3'd1 )+$signed( { 1'b0,x305 }  )+$signed( { 2'b0,x306 } <<<3'd1 )+$signed( -{ 1'b0,x308 } )+$signed( -{ 1'b0,x310 } )+$signed( -{ 3'b0,x311 }<<<3'd2)+$signed( -{ 1'b0,x312 } )+$signed( -{ 1'b0,x313 } )+$signed( -{ 3'b0,x314 }<<<3'd2)+$signed( { 2'b0,x315 } <<<3'd1 )+$signed( { 1'b0,x316 }  )+$signed( { 3'b0,x317 }<<<3'd2 )+$signed( { 4'b0,x318 }<<<3'd3 )+$signed( { 2'b0,x319 } <<<3'd1 )+$signed( { 2'b0,x321 } <<<3'd1 )+$signed( { 1'b0,x322 }  )+$signed( { 2'b0,x323 } <<<3'd1 )+$signed( -{ 1'b0,x324 } )+$signed( { 3'b0,x325 }<<<3'd2 )+$signed( { 2'b0,x327 } <<<3'd1 )+$signed( { 2'b0,x328 } <<<3'd1 )+$signed( -{ 1'b0,x329 } )+$signed( -{ 1'b0,x330 } )+$signed( -{ 2'b0,x331 }<<<3'd1 )+$signed( { 2'b0,x333 } <<<3'd1 )+$signed( { 1'b0,x334 }  )+$signed( -{ 2'b0,x335 }<<<3'd1 )+$signed( { 2'b0,x336 } <<<3'd1 )+$signed( { 1'b0,x337 }  )+$signed( { 1'b0,x338 }  )+$signed( -{ 2'b0,x339 }<<<3'd1 )+$signed( { 2'b0,x340 } <<<3'd1 )+$signed( { 1'b0,x341 }  )+$signed( -{ 3'b0,x342 }<<<3'd2)+$signed( { 3'b0,x343 }<<<3'd2 )+$signed( { 2'b0,x347 } <<<3'd1 )+$signed( { 3'b0,x348 }<<<3'd2 )+$signed( -{ 1'b0,x350 } )+$signed( { 1'b0,x351 }  )+$signed( -{ 2'b0,x352 }<<<3'd1 )+$signed( { 2'b0,x355 } <<<3'd1 )+$signed( { 3'b0,x356 }<<<3'd2 )+$signed( { 4'b0,x357 }<<<3'd3 )+$signed( { 3'b0,x358 }<<<3'd2 )+$signed( { 1'b0,x359 }  )+$signed( { 2'b0,x360 } <<<3'd1 )+$signed( { 1'b0,x361 }  )+$signed( -{ 3'b0,x362 }<<<3'd2)+$signed( -{ 3'b0,x363 }<<<3'd2)+$signed( -{ 2'b0,x364 }<<<3'd1 )+$signed( { 2'b0,x365 } <<<3'd1 )+$signed( { 1'b0,x366 }  )+$signed( -{ 1'b0,x367 } )+$signed( { 1'b0,x368 }  )+$signed( { 3'b0,x369 }<<<3'd2 )+$signed( { 3'b0,x370 }<<<3'd2 )+$signed( { 1'b0,x371 }  )+$signed( { 2'b0,x372 } <<<3'd1 )+$signed( { 2'b0,x374 } <<<3'd1 )+$signed( { 1'b0,x375 }  )+$signed( -{ 3'b0,x376 }<<<3'd2)+$signed( { 1'b0,x377 }  )+$signed( { 3'b0,x378 }<<<3'd2 )+$signed( { 3'b0,x379 }<<<3'd2 )+$signed( { 3'b0,x380 }<<<3'd2 )+$signed( { 2'b0,x381 } <<<3'd1 )+$signed( { 3'b0,x382 }<<<3'd2 )+$signed( { 3'b0,x383 }<<<3'd2 )+$signed( -{ 2'b0,x384 }<<<3'd1 )+$signed( { 2'b0,x385 } <<<3'd1 )+$signed( { 2'b0,x386 } <<<3'd1 )+$signed( { 3'b0,x388 }<<<3'd2 )+$signed( -{ 2'b0,x389 }<<<3'd1 )+$signed( { 3'b0,x390 }<<<3'd2 )+$signed( { 2'b0,x391 } <<<3'd1 )+$signed( -{ 2'b0,x392 }<<<3'd1 )+$signed( { 2'b0,x393 } <<<3'd1 )+$signed( -{ 1'b0,x394 } )+$signed( { 3'b0,x395 }<<<3'd2 )+$signed( -{ 2'b0,x396 }<<<3'd1 )+$signed( { 2'b0,x397 } <<<3'd1 )+$signed( -{ 2'b0,x398 }<<<3'd1 )+$signed( { 3'b0,x399 }<<<3'd2 )+$signed( { 2'b0,x400 } <<<3'd1 )+$signed( -{ 2'b0,x401 }<<<3'd1 )+$signed( { 1'b0,x403 }  )+$signed( -{ 3'b0,x404 }<<<3'd2)+$signed( { 3'b0,x406 }<<<3'd2 )+$signed( { 4'b0,x408 }<<<3'd3 )+$signed( { 1'b0,x409 }  )+$signed( { 2'b0,x410 } <<<3'd1 )+$signed( { 2'b0,x411 } <<<3'd1 )+$signed( { 2'b0,x412 } <<<3'd1 )+$signed( { 3'b0,x413 }<<<3'd2 )+$signed( { 3'b0,x414 }<<<3'd2 )+$signed( { 2'b0,x416 } <<<3'd1 )+$signed( -{ 2'b0,x417 }<<<3'd1 )+$signed( { 3'b0,x418 }<<<3'd2 )+$signed( { 3'b0,x419 }<<<3'd2 )+$signed( { 1'b0,x420 }  )+$signed( { 2'b0,x421 } <<<3'd1 )+$signed( { 1'b0,x423 }  )+$signed( { 2'b0,x425 } <<<3'd1 )+$signed( -{ 2'b0,x426 }<<<3'd1 )+$signed( { 2'b0,x427 } <<<3'd1 )+$signed( -{ 3'b0,x429 }<<<3'd2)+$signed( { 2'b0,x430 } <<<3'd1 )+$signed( { 3'b0,x431 }<<<3'd2 )+$signed( { 2'b0,x432 } <<<3'd1 )+$signed( -{ 2'b0,x434 }<<<3'd1 )+$signed( -{ 3'b0,x435 }<<<3'd2)+$signed( { 1'b0,x436 }  )+$signed( -{ 1'b0,x437 } )+$signed( { 2'b0,x438 } <<<3'd1 )+$signed( -{ 2'b0,x439 }<<<3'd1 )+$signed( { 2'b0,x440 } <<<3'd1 )+$signed( { 2'b0,x441 } <<<3'd1 )+$signed( { 2'b0,x442 } <<<3'd1 )+$signed( { 1'b0,x443 }  )+$signed( { 3'b0,x444 }<<<3'd2 )+$signed( -{ 2'b0,x445 }<<<3'd1 )+$signed( { 1'b0,x447 }  )+$signed( { 1'b0,x448 }  )+$signed( -{ 2'b0,x449 }<<<3'd1 )+$signed( -{ 1'b0,x450 } )+$signed( { 4'b0,x452 }<<<3'd3 )+$signed( -{ 2'b0,x453 }<<<3'd1 )+$signed( -{ 3'b0,x454 }<<<3'd2)+$signed( { 4'b0,x455 }<<<3'd3 )+$signed( -{ 1'b0,x456 } )+$signed( { 3'b0,x457 }<<<3'd2 )+$signed( { 2'b0,x459 } <<<3'd1 )+$signed( -{ 1'b0,x460 } )+$signed( -{ 2'b0,x461 }<<<3'd1 )+$signed( { 3'b0,x463 }<<<3'd2 )+$signed( { 2'b0,x464 } <<<3'd1 )+$signed( { 4'b0,x465 }<<<3'd3 )+$signed( { 2'b0,x467 } <<<3'd1 )+$signed( -{ 1'b0,x468 } )+$signed( { 1'b0,x469 }  )+$signed( { 2'b0,x471 } <<<3'd1 )+$signed( { 3'b0,x472 }<<<3'd2 )+$signed( { 1'b0,x473 }  )+$signed( -{ 1'b0,x474 } )+$signed( { 1'b0,x476 }  )+$signed( { 3'b0,x477 }<<<3'd2 )+$signed( -{ 1'b0,x478 } )+$signed( -{ 1'b0,x479 } )+$signed( { 3'b0,x480 }<<<3'd2 )+$signed( { 2'b0,x481 } <<<3'd1 )+$signed( { 2'b0,x482 } <<<3'd1 )+$signed( { 3'b0,x483 }<<<3'd2 )+$signed( { 2'b0,x484 } <<<3'd1 )+$signed( -{ 1'b0,x486 } )+$signed( { 2'b0,x487 } <<<3'd1 )+$signed( { 1'b0,x488 }  )+$signed( -{ 3'b0,x489 }<<<3'd2)+$signed( { 3'b0,x490 }<<<3'd2 )+$signed( -{ 2'b0,x491 }<<<3'd1 )+$signed( { 2'b0,x492 } <<<3'd1 )+$signed( { 1'b0,x493 }  )+$signed( { 3'b0,x494 }<<<3'd2 )+$signed( -{ 4'b0, x495 }<<<3'd3 )-$signed(13'd48);
assign y11=temp_y[11][13] ==1'b1 ? 6'd0 :  
    temp_y[11][10] ==1'b1 ? 6'd63 : 
    temp_y[11][3]==1'b1 ? temp_y[11][9:4]+1'b1 : temp_y[11][9:4];
assign temp_y[12] = 
+$signed( { 1'b0,x0 }  )+$signed( -{ 2'b0,x1 }<<<3'd1 )+$signed( { 1'b0,x3 }  )+$signed( -{ 1'b0,x4 } )+$signed( -{ 2'b0,x5 }<<<3'd1 )+$signed( -{ 1'b0,x6 } )+$signed( { 3'b0,x7 }<<<3'd2 )+$signed( { 1'b0,x8 }  )+$signed( -{ 1'b0,x9 } )+$signed( { 3'b0,x10 }<<<3'd2 )+$signed( { 1'b0,x11 }  )+$signed( -{ 2'b0,x12 }<<<3'd1 )+$signed( -{ 2'b0,x13 }<<<3'd1 )+$signed( -{ 2'b0,x14 }<<<3'd1 )+$signed( { 3'b0,x15 }<<<3'd2 )+$signed( { 1'b0,x16 }  )+$signed( { 2'b0,x18 } <<<3'd1 )+$signed( { 1'b0,x19 }  )+$signed( -{ 1'b0,x20 } )+$signed( { 1'b0,x21 }  )+$signed( { 3'b0,x22 }<<<3'd2 )+$signed( { 1'b0,x23 }  )+$signed( { 1'b0,x25 }  )+$signed( { 1'b0,x26 }  )+$signed( -{ 2'b0,x27 }<<<3'd1 )+$signed( -{ 3'b0,x28 }<<<3'd2)+$signed( { 2'b0,x29 } <<<3'd1 )+$signed( -{ 1'b0,x30 } )+$signed( { 2'b0,x31 } <<<3'd1 )+$signed( { 2'b0,x32 } <<<3'd1 )+$signed( { 2'b0,x33 } <<<3'd1 )+$signed( { 3'b0,x34 }<<<3'd2 )+$signed( { 1'b0,x35 }  )+$signed( { 1'b0,x38 }  )+$signed( { 2'b0,x39 } <<<3'd1 )+$signed( { 1'b0,x40 }  )+$signed( { 1'b0,x42 }  )+$signed( { 3'b0,x43 }<<<3'd2 )+$signed( { 1'b0,x45 }  )+$signed( { 1'b0,x46 }  )+$signed( { 2'b0,x47 } <<<3'd1 )+$signed( { 2'b0,x49 } <<<3'd1 )+$signed( { 1'b0,x50 }  )+$signed( { 3'b0,x51 }<<<3'd2 )+$signed( { 1'b0,x53 }  )+$signed( { 3'b0,x54 }<<<3'd2 )+$signed( -{ 2'b0,x55 }<<<3'd1 )+$signed( { 1'b0,x56 }  )+$signed( { 1'b0,x57 }  )+$signed( { 1'b0,x58 }  )+$signed( -{ 2'b0,x59 }<<<3'd1 )+$signed( -{ 1'b0,x60 } )+$signed( { 2'b0,x61 } <<<3'd1 )+$signed( { 2'b0,x62 } <<<3'd1 )+$signed( { 1'b0,x63 }  )+$signed( { 1'b0,x64 }  )+$signed( { 1'b0,x65 }  )+$signed( -{ 1'b0,x67 } )+$signed( -{ 2'b0,x68 }<<<3'd1 )+$signed( { 1'b0,x71 }  )+$signed( -{ 1'b0,x73 } )+$signed( { 3'b0,x74 }<<<3'd2 )+$signed( { 1'b0,x75 }  )+$signed( { 3'b0,x76 }<<<3'd2 )+$signed( -{ 1'b0,x78 } )+$signed( -{ 2'b0,x79 }<<<3'd1 )+$signed( { 1'b0,x80 }  )+$signed( { 1'b0,x81 }  )+$signed( { 2'b0,x83 } <<<3'd1 )+$signed( -{ 3'b0,x84 }<<<3'd2)+$signed( -{ 2'b0,x85 }<<<3'd1 )+$signed( { 3'b0,x87 }<<<3'd2 )+$signed( -{ 1'b0,x89 } )+$signed( -{ 3'b0,x91 }<<<3'd2)+$signed( { 3'b0,x92 }<<<3'd2 )+$signed( -{ 3'b0,x93 }<<<3'd2)+$signed( { 3'b0,x94 }<<<3'd2 )+$signed( { 3'b0,x95 }<<<3'd2 )+$signed( { 3'b0,x96 }<<<3'd2 )+$signed( { 4'b0,x97 }<<<3'd3 )+$signed( -{ 2'b0,x98 }<<<3'd1 )+$signed( -{ 3'b0,x99 }<<<3'd2)+$signed( -{ 4'b0, x100 }<<<3'd3 )+$signed( { 3'b0,x101 }<<<3'd2 )+$signed( -{ 3'b0,x102 }<<<3'd2)+$signed( -{ 2'b0,x103 }<<<3'd1 )+$signed( { 1'b0,x104 }  )+$signed( { 2'b0,x105 } <<<3'd1 )+$signed( { 3'b0,x106 }<<<3'd2 )+$signed( { 1'b0,x108 }  )+$signed( { 3'b0,x110 }<<<3'd2 )+$signed( -{ 2'b0,x111 }<<<3'd1 )+$signed( { 1'b0,x112 }  )+$signed( { 2'b0,x113 } <<<3'd1 )+$signed( { 3'b0,x114 }<<<3'd2 )+$signed( { 4'b0,x115 }<<<3'd3 )+$signed( -{ 1'b0,x116 } )+$signed( -{ 3'b0,x117 }<<<3'd2)+$signed( -{ 4'b0, x118 }<<<3'd3 )+$signed( { 3'b0,x119 }<<<3'd2 )+$signed( -{ 3'b0,x120 }<<<3'd2)+$signed( -{ 2'b0,x121 }<<<3'd1 )+$signed( { 1'b0,x122 }  )+$signed( { 3'b0,x123 }<<<3'd2 )+$signed( -{ 2'b0,x124 }<<<3'd1 )+$signed( { 2'b0,x125 } <<<3'd1 )+$signed( -{ 2'b0,x126 }<<<3'd1 )+$signed( -{ 1'b0,x127 } )+$signed( { 2'b0,x128 } <<<3'd1 )+$signed( { 1'b0,x130 }  )+$signed( -{ 1'b0,x131 } )+$signed( { 3'b0,x133 }<<<3'd2 )+$signed( { 1'b0,x134 }  )+$signed( { 1'b0,x135 }  )+$signed( -{ 2'b0,x137 }<<<3'd1 )+$signed( -{ 2'b0,x138 }<<<3'd1 )+$signed( { 1'b0,x139 }  )+$signed( { 1'b0,x140 }  )+$signed( { 2'b0,x141 } <<<3'd1 )+$signed( { 3'b0,x143 }<<<3'd2 )+$signed( { 1'b0,x145 }  )+$signed( { 3'b0,x146 }<<<3'd2 )+$signed( { 2'b0,x147 } <<<3'd1 )+$signed( { 2'b0,x148 } <<<3'd1 )+$signed( { 1'b0,x149 }  )+$signed( { 2'b0,x151 } <<<3'd1 )+$signed( { 1'b0,x152 }  )+$signed( { 2'b0,x153 } <<<3'd1 )+$signed( { 3'b0,x154 }<<<3'd2 )+$signed( { 1'b0,x155 }  )+$signed( { 1'b0,x156 }  )+$signed( -{ 1'b0,x157 } )+$signed( { 2'b0,x159 } <<<3'd1 )+$signed( -{ 3'b0,x160 }<<<3'd2)+$signed( { 2'b0,x161 } <<<3'd1 )+$signed( -{ 1'b0,x162 } )+$signed( -{ 3'b0,x163 }<<<3'd2)+$signed( { 2'b0,x164 } <<<3'd1 )+$signed( -{ 2'b0,x165 }<<<3'd1 )+$signed( { 3'b0,x166 }<<<3'd2 )+$signed( { 3'b0,x167 }<<<3'd2 )+$signed( { 3'b0,x168 }<<<3'd2 )+$signed( -{ 2'b0,x170 }<<<3'd1 )+$signed( -{ 3'b0,x171 }<<<3'd2)+$signed( { 4'b0,x173 }<<<3'd3 )+$signed( -{ 3'b0,x174 }<<<3'd2)+$signed( -{ 3'b0,x175 }<<<3'd2)+$signed( -{ 3'b0,x176 }<<<3'd2)+$signed( { 3'b0,x177 }<<<3'd2 )+$signed( -{ 3'b0,x178 }<<<3'd2)+$signed( { 2'b0,x179 } <<<3'd1 )+$signed( -{ 2'b0,x181 }<<<3'd1 )+$signed( { 2'b0,x182 } <<<3'd1 )+$signed( { 2'b0,x183 } <<<3'd1 )+$signed( -{ 2'b0,x184 }<<<3'd1 )+$signed( { 2'b0,x185 } <<<3'd1 )+$signed( { 2'b0,x186 } <<<3'd1 )+$signed( { 2'b0,x187 } <<<3'd1 )+$signed( -{ 4'b0, x189 }<<<3'd3 )+$signed( { 3'b0,x191 }<<<3'd2 )+$signed( -{ 3'b0,x192 }<<<3'd2)+$signed( -{ 2'b0,x193 }<<<3'd1 )+$signed( -{ 3'b0,x194 }<<<3'd2)+$signed( { 2'b0,x195 } <<<3'd1 )+$signed( { 2'b0,x196 } <<<3'd1 )+$signed( { 2'b0,x197 } <<<3'd1 )+$signed( { 2'b0,x198 } <<<3'd1 )+$signed( -{ 3'b0,x199 }<<<3'd2)+$signed( { 2'b0,x201 } <<<3'd1 )+$signed( { 2'b0,x202 } <<<3'd1 )+$signed( { 1'b0,x204 }  )+$signed( { 1'b0,x205 }  )+$signed( { 1'b0,x206 }  )+$signed( -{ 1'b0,x207 } )+$signed( -{ 1'b0,x209 } )+$signed( -{ 2'b0,x210 }<<<3'd1 )+$signed( -{ 2'b0,x211 }<<<3'd1 )+$signed( { 2'b0,x213 } <<<3'd1 )+$signed( { 2'b0,x214 } <<<3'd1 )+$signed( { 3'b0,x215 }<<<3'd2 )+$signed( { 2'b0,x216 } <<<3'd1 )+$signed( { 3'b0,x217 }<<<3'd2 )+$signed( { 3'b0,x218 }<<<3'd2 )+$signed( -{ 1'b0,x219 } )+$signed( { 3'b0,x220 }<<<3'd2 )+$signed( -{ 3'b0,x222 }<<<3'd2)+$signed( { 2'b0,x223 } <<<3'd1 )+$signed( -{ 1'b0,x224 } )+$signed( { 3'b0,x225 }<<<3'd2 )+$signed( { 2'b0,x226 } <<<3'd1 )+$signed( { 2'b0,x227 } <<<3'd1 )+$signed( -{ 1'b0,x228 } )+$signed( -{ 2'b0,x230 }<<<3'd1 )+$signed( { 3'b0,x231 }<<<3'd2 )+$signed( -{ 1'b0,x232 } )+$signed( { 2'b0,x234 } <<<3'd1 )+$signed( -{ 2'b0,x235 }<<<3'd1 )+$signed( { 2'b0,x236 } <<<3'd1 )+$signed( -{ 2'b0,x237 }<<<3'd1 )+$signed( { 4'b0,x238 }<<<3'd3 )+$signed( { 2'b0,x239 } <<<3'd1 )+$signed( { 3'b0,x240 }<<<3'd2 )+$signed( -{ 3'b0,x241 }<<<3'd2)+$signed( { 1'b0,x244 }  )+$signed( { 3'b0,x245 }<<<3'd2 )+$signed( -{ 1'b0,x246 } )+$signed( { 2'b0,x247 } <<<3'd1 )+$signed( -{ 2'b0,x248 }<<<3'd1 )+$signed( { 2'b0,x249 } <<<3'd1 )+$signed( { 1'b0,x251 }  )+$signed( { 2'b0,x254 } <<<3'd1 )+$signed( -{ 1'b0,x256 } )+$signed( { 1'b0,x257 }  )+$signed( { 2'b0,x258 } <<<3'd1 )+$signed( -{ 3'b0,x259 }<<<3'd2)+$signed( { 2'b0,x260 } <<<3'd1 )+$signed( -{ 2'b0,x261 }<<<3'd1 )+$signed( { 1'b0,x262 }  )+$signed( { 2'b0,x263 } <<<3'd1 )+$signed( -{ 2'b0,x264 }<<<3'd1 )+$signed( { 3'b0,x265 }<<<3'd2 )+$signed( -{ 2'b0,x266 }<<<3'd1 )+$signed( { 1'b0,x267 }  )+$signed( -{ 2'b0,x268 }<<<3'd1 )+$signed( { 2'b0,x269 } <<<3'd1 )+$signed( { 2'b0,x270 } <<<3'd1 )+$signed( { 1'b0,x271 }  )+$signed( -{ 1'b0,x272 } )+$signed( -{ 1'b0,x273 } )+$signed( { 2'b0,x274 } <<<3'd1 )+$signed( -{ 2'b0,x275 }<<<3'd1 )+$signed( -{ 1'b0,x276 } )+$signed( -{ 2'b0,x277 }<<<3'd1 )+$signed( { 2'b0,x279 } <<<3'd1 )+$signed( { 2'b0,x280 } <<<3'd1 )+$signed( -{ 1'b0,x281 } )+$signed( { 2'b0,x282 } <<<3'd1 )+$signed( -{ 2'b0,x284 }<<<3'd1 )+$signed( { 2'b0,x285 } <<<3'd1 )+$signed( -{ 1'b0,x286 } )+$signed( { 2'b0,x287 } <<<3'd1 )+$signed( { 2'b0,x288 } <<<3'd1 )+$signed( { 1'b0,x289 }  )+$signed( { 2'b0,x290 } <<<3'd1 )+$signed( { 1'b0,x291 }  )+$signed( -{ 1'b0,x292 } )+$signed( -{ 1'b0,x293 } )+$signed( { 1'b0,x294 }  )+$signed( { 3'b0,x296 }<<<3'd2 )+$signed( { 1'b0,x298 }  )+$signed( { 2'b0,x299 } <<<3'd1 )+$signed( { 1'b0,x300 }  )+$signed( { 3'b0,x301 }<<<3'd2 )+$signed( -{ 1'b0,x302 } )+$signed( { 1'b0,x303 }  )+$signed( { 2'b0,x304 } <<<3'd1 )+$signed( { 3'b0,x305 }<<<3'd2 )+$signed( -{ 1'b0,x306 } )+$signed( { 3'b0,x307 }<<<3'd2 )+$signed( { 2'b0,x308 } <<<3'd1 )+$signed( { 3'b0,x309 }<<<3'd2 )+$signed( -{ 2'b0,x310 }<<<3'd1 )+$signed( { 3'b0,x311 }<<<3'd2 )+$signed( { 1'b0,x312 }  )+$signed( { 1'b0,x313 }  )+$signed( -{ 2'b0,x315 }<<<3'd1 )+$signed( { 2'b0,x316 } <<<3'd1 )+$signed( { 3'b0,x317 }<<<3'd2 )+$signed( { 3'b0,x318 }<<<3'd2 )+$signed( { 1'b0,x320 }  )+$signed( -{ 2'b0,x321 }<<<3'd1 )+$signed( { 1'b0,x322 }  )+$signed( -{ 2'b0,x323 }<<<3'd1 )+$signed( { 2'b0,x326 } <<<3'd1 )+$signed( -{ 1'b0,x328 } )+$signed( { 2'b0,x330 } <<<3'd1 )+$signed( { 3'b0,x331 }<<<3'd2 )+$signed( -{ 3'b0,x332 }<<<3'd2)+$signed( { 2'b0,x333 } <<<3'd1 )+$signed( { 1'b0,x336 }  )+$signed( -{ 1'b0,x337 } )+$signed( { 1'b0,x338 }  )+$signed( { 1'b0,x340 }  )+$signed( -{ 1'b0,x341 } )+$signed( { 2'b0,x342 } <<<3'd1 )+$signed( { 1'b0,x343 }  )+$signed( -{ 1'b0,x344 } )+$signed( -{ 2'b0,x345 }<<<3'd1 )+$signed( { 3'b0,x346 }<<<3'd2 )+$signed( { 1'b0,x347 }  )+$signed( { 1'b0,x348 }  )+$signed( { 2'b0,x349 } <<<3'd1 )+$signed( { 1'b0,x350 }  )+$signed( -{ 2'b0,x351 }<<<3'd1 )+$signed( { 2'b0,x352 } <<<3'd1 )+$signed( -{ 3'b0,x353 }<<<3'd2)+$signed( { 2'b0,x354 } <<<3'd1 )+$signed( -{ 1'b0,x357 } )+$signed( -{ 1'b0,x358 } )+$signed( { 3'b0,x359 }<<<3'd2 )+$signed( { 1'b0,x360 }  )+$signed( { 3'b0,x361 }<<<3'd2 )+$signed( -{ 4'b0, x362 }<<<3'd3 )+$signed( { 1'b0,x363 }  )+$signed( { 3'b0,x364 }<<<3'd2 )+$signed( { 2'b0,x365 } <<<3'd1 )+$signed( -{ 1'b0,x366 } )+$signed( { 1'b0,x367 }  )+$signed( { 1'b0,x369 }  )+$signed( { 4'b0,x370 }<<<3'd3 )+$signed( { 1'b0,x371 }  )+$signed( { 2'b0,x372 } <<<3'd1 )+$signed( { 2'b0,x374 } <<<3'd1 )+$signed( -{ 3'b0,x375 }<<<3'd2)+$signed( { 3'b0,x376 }<<<3'd2 )+$signed( { 3'b0,x377 }<<<3'd2 )+$signed( { 3'b0,x378 }<<<3'd2 )+$signed( -{ 2'b0,x379 }<<<3'd1 )+$signed( { 2'b0,x381 } <<<3'd1 )+$signed( { 1'b0,x382 }  )+$signed( { 2'b0,x383 } <<<3'd1 )+$signed( -{ 1'b0,x384 } )+$signed( { 3'b0,x385 }<<<3'd2 )+$signed( -{ 3'b0,x386 }<<<3'd2)+$signed( { 3'b0,x387 }<<<3'd2 )+$signed( { 2'b0,x388 } <<<3'd1 )+$signed( { 2'b0,x389 } <<<3'd1 )+$signed( { 1'b0,x390 }  )+$signed( { 2'b0,x392 } <<<3'd1 )+$signed( -{ 3'b0,x393 }<<<3'd2)+$signed( { 3'b0,x394 }<<<3'd2 )+$signed( -{ 1'b0,x395 } )+$signed( -{ 2'b0,x396 }<<<3'd1 )+$signed( -{ 2'b0,x397 }<<<3'd1 )+$signed( { 2'b0,x398 } <<<3'd1 )+$signed( -{ 2'b0,x399 }<<<3'd1 )+$signed( { 1'b0,x401 }  )+$signed( { 1'b0,x402 }  )+$signed( { 2'b0,x403 } <<<3'd1 )+$signed( { 3'b0,x404 }<<<3'd2 )+$signed( -{ 2'b0,x405 }<<<3'd1 )+$signed( -{ 3'b0,x406 }<<<3'd2)+$signed( { 2'b0,x407 } <<<3'd1 )+$signed( { 1'b0,x408 }  )+$signed( -{ 3'b0,x410 }<<<3'd2)+$signed( { 2'b0,x411 } <<<3'd1 )+$signed( -{ 2'b0,x412 }<<<3'd1 )+$signed( -{ 2'b0,x413 }<<<3'd1 )+$signed( -{ 3'b0,x414 }<<<3'd2)+$signed( { 3'b0,x415 }<<<3'd2 )+$signed( { 2'b0,x416 } <<<3'd1 )+$signed( { 3'b0,x417 }<<<3'd2 )+$signed( -{ 1'b0,x418 } )+$signed( -{ 2'b0,x419 }<<<3'd1 )+$signed( { 2'b0,x420 } <<<3'd1 )+$signed( { 3'b0,x422 }<<<3'd2 )+$signed( -{ 2'b0,x423 }<<<3'd1 )+$signed( { 3'b0,x424 }<<<3'd2 )+$signed( -{ 2'b0,x425 }<<<3'd1 )+$signed( -{ 2'b0,x426 }<<<3'd1 )+$signed( -{ 1'b0,x427 } )+$signed( { 1'b0,x428 }  )+$signed( { 3'b0,x429 }<<<3'd2 )+$signed( { 3'b0,x430 }<<<3'd2 )+$signed( -{ 3'b0,x431 }<<<3'd2)+$signed( { 2'b0,x433 } <<<3'd1 )+$signed( { 2'b0,x434 } <<<3'd1 )+$signed( { 3'b0,x435 }<<<3'd2 )+$signed( -{ 3'b0,x436 }<<<3'd2)+$signed( { 1'b0,x437 }  )+$signed( -{ 3'b0,x438 }<<<3'd2)+$signed( { 3'b0,x439 }<<<3'd2 )+$signed( { 2'b0,x441 } <<<3'd1 )+$signed( { 3'b0,x443 }<<<3'd2 )+$signed( { 3'b0,x444 }<<<3'd2 )+$signed( { 1'b0,x446 }  )+$signed( -{ 2'b0,x447 }<<<3'd1 )+$signed( -{ 2'b0,x448 }<<<3'd1 )+$signed( { 1'b0,x450 }  )+$signed( -{ 1'b0,x451 } )+$signed( -{ 2'b0,x452 }<<<3'd1 )+$signed( { 1'b0,x454 }  )+$signed( -{ 3'b0,x455 }<<<3'd2)+$signed( { 2'b0,x456 } <<<3'd1 )+$signed( -{ 3'b0,x457 }<<<3'd2)+$signed( -{ 2'b0,x458 }<<<3'd1 )+$signed( { 2'b0,x459 } <<<3'd1 )+$signed( -{ 1'b0,x460 } )+$signed( { 2'b0,x461 } <<<3'd1 )+$signed( -{ 1'b0,x462 } )+$signed( { 1'b0,x463 }  )+$signed( -{ 3'b0,x464 }<<<3'd2)+$signed( -{ 2'b0,x465 }<<<3'd1 )+$signed( { 2'b0,x466 } <<<3'd1 )+$signed( { 2'b0,x467 } <<<3'd1 )+$signed( { 1'b0,x468 }  )+$signed( -{ 2'b0,x469 }<<<3'd1 )+$signed( -{ 2'b0,x470 }<<<3'd1 )+$signed( { 2'b0,x471 } <<<3'd1 )+$signed( -{ 1'b0,x473 } )+$signed( -{ 2'b0,x474 }<<<3'd1 )+$signed( { 2'b0,x475 } <<<3'd1 )+$signed( { 3'b0,x476 }<<<3'd2 )+$signed( -{ 1'b0,x477 } )+$signed( { 2'b0,x479 } <<<3'd1 )+$signed( { 1'b0,x480 }  )+$signed( -{ 2'b0,x481 }<<<3'd1 )+$signed( { 3'b0,x482 }<<<3'd2 )+$signed( -{ 2'b0,x483 }<<<3'd1 )+$signed( -{ 3'b0,x484 }<<<3'd2)+$signed( -{ 2'b0,x485 }<<<3'd1 )+$signed( { 2'b0,x486 } <<<3'd1 )+$signed( { 3'b0,x487 }<<<3'd2 )+$signed( -{ 3'b0,x488 }<<<3'd2)+$signed( { 3'b0,x489 }<<<3'd2 )+$signed( -{ 2'b0,x490 }<<<3'd1 )+$signed( { 2'b0,x491 } <<<3'd1 )+$signed( { 1'b0,x492 }  )+$signed( { 2'b0,x493 } <<<3'd1 )+$signed( -{ 1'b0,x494 } )+$signed( { 4'b0,x495 }<<<3'd3 )-$signed(13'd8);
assign y12=temp_y[12][13] ==1'b1 ? 6'd0 :  
    temp_y[12][10] ==1'b1 ? 6'd63 : 
    temp_y[12][3]==1'b1 ? temp_y[12][9:4]+1'b1 : temp_y[12][9:4];
assign temp_y[13] = 
+$signed( -{ 2'b0,x0 }<<<3'd1 )+$signed( { 2'b0,x1 } <<<3'd1 )+$signed( -{ 2'b0,x2 }<<<3'd1 )+$signed( -{ 2'b0,x3 }<<<3'd1 )+$signed( -{ 2'b0,x4 }<<<3'd1 )+$signed( -{ 1'b0,x5 } )+$signed( -{ 2'b0,x6 }<<<3'd1 )+$signed( -{ 2'b0,x7 }<<<3'd1 )+$signed( -{ 1'b0,x8 } )+$signed( -{ 2'b0,x9 }<<<3'd1 )+$signed( -{ 2'b0,x10 }<<<3'd1 )+$signed( { 3'b0,x11 }<<<3'd2 )+$signed( -{ 1'b0,x12 } )+$signed( { 2'b0,x13 } <<<3'd1 )+$signed( { 3'b0,x14 }<<<3'd2 )+$signed( { 3'b0,x15 }<<<3'd2 )+$signed( -{ 2'b0,x16 }<<<3'd1 )+$signed( { 1'b0,x17 }  )+$signed( -{ 2'b0,x18 }<<<3'd1 )+$signed( { 3'b0,x19 }<<<3'd2 )+$signed( -{ 1'b0,x20 } )+$signed( { 2'b0,x21 } <<<3'd1 )+$signed( { 2'b0,x22 } <<<3'd1 )+$signed( -{ 2'b0,x23 }<<<3'd1 )+$signed( -{ 4'b0, x25 }<<<3'd3 )+$signed( -{ 3'b0,x27 }<<<3'd2)+$signed( { 3'b0,x28 }<<<3'd2 )+$signed( { 3'b0,x29 }<<<3'd2 )+$signed( -{ 2'b0,x31 }<<<3'd1 )+$signed( -{ 1'b0,x35 } )+$signed( -{ 2'b0,x36 }<<<3'd1 )+$signed( { 3'b0,x37 }<<<3'd2 )+$signed( -{ 2'b0,x39 }<<<3'd1 )+$signed( -{ 1'b0,x41 } )+$signed( { 1'b0,x42 }  )+$signed( { 1'b0,x43 }  )+$signed( -{ 1'b0,x44 } )+$signed( -{ 3'b0,x45 }<<<3'd2)+$signed( { 3'b0,x46 }<<<3'd2 )+$signed( { 3'b0,x47 }<<<3'd2 )+$signed( { 2'b0,x48 } <<<3'd1 )+$signed( -{ 2'b0,x49 }<<<3'd1 )+$signed( { 2'b0,x50 } <<<3'd1 )+$signed( { 3'b0,x51 }<<<3'd2 )+$signed( -{ 3'b0,x52 }<<<3'd2)+$signed( { 1'b0,x53 }  )+$signed( { 3'b0,x54 }<<<3'd2 )+$signed( { 3'b0,x55 }<<<3'd2 )+$signed( { 2'b0,x56 } <<<3'd1 )+$signed( -{ 2'b0,x57 }<<<3'd1 )+$signed( { 2'b0,x58 } <<<3'd1 )+$signed( -{ 2'b0,x59 }<<<3'd1 )+$signed( { 1'b0,x60 }  )+$signed( -{ 1'b0,x61 } )+$signed( -{ 1'b0,x62 } )+$signed( { 1'b0,x63 }  )+$signed( -{ 2'b0,x64 }<<<3'd1 )+$signed( { 3'b0,x65 }<<<3'd2 )+$signed( { 3'b0,x66 }<<<3'd2 )+$signed( { 1'b0,x68 }  )+$signed( { 3'b0,x69 }<<<3'd2 )+$signed( { 3'b0,x70 }<<<3'd2 )+$signed( { 2'b0,x71 } <<<3'd1 )+$signed( { 2'b0,x72 } <<<3'd1 )+$signed( { 2'b0,x73 } <<<3'd1 )+$signed( -{ 3'b0,x74 }<<<3'd2)+$signed( { 3'b0,x75 }<<<3'd2 )+$signed( -{ 3'b0,x76 }<<<3'd2)+$signed( { 1'b0,x77 }  )+$signed( { 3'b0,x78 }<<<3'd2 )+$signed( -{ 3'b0,x79 }<<<3'd2)+$signed( { 1'b0,x81 }  )+$signed( -{ 1'b0,x82 } )+$signed( { 2'b0,x83 } <<<3'd1 )+$signed( { 3'b0,x84 }<<<3'd2 )+$signed( { 1'b0,x85 }  )+$signed( { 1'b0,x86 }  )+$signed( { 1'b0,x87 }  )+$signed( { 3'b0,x88 }<<<3'd2 )+$signed( { 2'b0,x89 } <<<3'd1 )+$signed( { 2'b0,x91 } <<<3'd1 )+$signed( -{ 1'b0,x92 } )+$signed( -{ 2'b0,x93 }<<<3'd1 )+$signed( { 2'b0,x94 } <<<3'd1 )+$signed( -{ 3'b0,x95 }<<<3'd2)+$signed( { 2'b0,x96 } <<<3'd1 )+$signed( -{ 2'b0,x97 }<<<3'd1 )+$signed( { 3'b0,x98 }<<<3'd2 )+$signed( -{ 3'b0,x99 }<<<3'd2)+$signed( { 1'b0,x100 }  )+$signed( { 1'b0,x101 }  )+$signed( { 2'b0,x102 } <<<3'd1 )+$signed( { 2'b0,x103 } <<<3'd1 )+$signed( { 2'b0,x104 } <<<3'd1 )+$signed( -{ 2'b0,x105 }<<<3'd1 )+$signed( -{ 2'b0,x106 }<<<3'd1 )+$signed( { 2'b0,x107 } <<<3'd1 )+$signed( { 2'b0,x108 } <<<3'd1 )+$signed( { 2'b0,x109 } <<<3'd1 )+$signed( { 1'b0,x111 }  )+$signed( -{ 2'b0,x112 }<<<3'd1 )+$signed( -{ 3'b0,x113 }<<<3'd2)+$signed( -{ 3'b0,x114 }<<<3'd2)+$signed( -{ 4'b0, x115 }<<<3'd3 )+$signed( -{ 2'b0,x117 }<<<3'd1 )+$signed( { 4'b0,x118 }<<<3'd3 )+$signed( { 2'b0,x119 } <<<3'd1 )+$signed( { 3'b0,x120 }<<<3'd2 )+$signed( { 2'b0,x121 } <<<3'd1 )+$signed( { 2'b0,x122 } <<<3'd1 )+$signed( { 1'b0,x123 }  )+$signed( -{ 2'b0,x124 }<<<3'd1 )+$signed( { 2'b0,x125 } <<<3'd1 )+$signed( -{ 1'b0,x126 } )+$signed( { 2'b0,x127 } <<<3'd1 )+$signed( { 1'b0,x128 }  )+$signed( -{ 1'b0,x129 } )+$signed( -{ 3'b0,x130 }<<<3'd2)+$signed( -{ 1'b0,x131 } )+$signed( -{ 1'b0,x132 } )+$signed( -{ 2'b0,x133 }<<<3'd1 )+$signed( -{ 1'b0,x134 } )+$signed( { 1'b0,x135 }  )+$signed( { 1'b0,x136 }  )+$signed( { 2'b0,x137 } <<<3'd1 )+$signed( { 3'b0,x138 }<<<3'd2 )+$signed( { 3'b0,x139 }<<<3'd2 )+$signed( { 1'b0,x142 }  )+$signed( { 1'b0,x143 }  )+$signed( -{ 3'b0,x144 }<<<3'd2)+$signed( { 3'b0,x145 }<<<3'd2 )+$signed( { 1'b0,x146 }  )+$signed( { 1'b0,x147 }  )+$signed( -{ 2'b0,x148 }<<<3'd1 )+$signed( { 2'b0,x149 } <<<3'd1 )+$signed( -{ 1'b0,x150 } )+$signed( -{ 1'b0,x151 } )+$signed( -{ 3'b0,x152 }<<<3'd2)+$signed( { 2'b0,x153 } <<<3'd1 )+$signed( { 2'b0,x154 } <<<3'd1 )+$signed( { 1'b0,x155 }  )+$signed( { 3'b0,x156 }<<<3'd2 )+$signed( { 1'b0,x158 }  )+$signed( -{ 1'b0,x159 } )+$signed( { 3'b0,x160 }<<<3'd2 )+$signed( { 3'b0,x163 }<<<3'd2 )+$signed( { 1'b0,x164 }  )+$signed( { 2'b0,x165 } <<<3'd1 )+$signed( -{ 2'b0,x166 }<<<3'd1 )+$signed( { 2'b0,x167 } <<<3'd1 )+$signed( -{ 1'b0,x168 } )+$signed( -{ 1'b0,x169 } )+$signed( -{ 3'b0,x170 }<<<3'd2)+$signed( { 1'b0,x171 }  )+$signed( { 3'b0,x172 }<<<3'd2 )+$signed( { 3'b0,x173 }<<<3'd2 )+$signed( { 3'b0,x174 }<<<3'd2 )+$signed( { 2'b0,x175 } <<<3'd1 )+$signed( { 1'b0,x176 }  )+$signed( -{ 1'b0,x177 } )+$signed( -{ 1'b0,x178 } )+$signed( -{ 1'b0,x179 } )+$signed( -{ 3'b0,x182 }<<<3'd2)+$signed( { 3'b0,x183 }<<<3'd2 )+$signed( -{ 2'b0,x184 }<<<3'd1 )+$signed( { 2'b0,x185 } <<<3'd1 )+$signed( -{ 3'b0,x186 }<<<3'd2)+$signed( -{ 2'b0,x187 }<<<3'd1 )+$signed( -{ 3'b0,x188 }<<<3'd2)+$signed( { 2'b0,x189 } <<<3'd1 )+$signed( { 3'b0,x190 }<<<3'd2 )+$signed( { 3'b0,x191 }<<<3'd2 )+$signed( { 3'b0,x192 }<<<3'd2 )+$signed( { 2'b0,x193 } <<<3'd1 )+$signed( -{ 2'b0,x195 }<<<3'd1 )+$signed( { 3'b0,x196 }<<<3'd2 )+$signed( { 1'b0,x198 }  )+$signed( { 3'b0,x199 }<<<3'd2 )+$signed( { 2'b0,x200 } <<<3'd1 )+$signed( -{ 2'b0,x201 }<<<3'd1 )+$signed( { 2'b0,x202 } <<<3'd1 )+$signed( { 2'b0,x205 } <<<3'd1 )+$signed( -{ 3'b0,x206 }<<<3'd2)+$signed( { 3'b0,x208 }<<<3'd2 )+$signed( { 2'b0,x209 } <<<3'd1 )+$signed( { 3'b0,x210 }<<<3'd2 )+$signed( { 2'b0,x211 } <<<3'd1 )+$signed( { 2'b0,x212 } <<<3'd1 )+$signed( { 1'b0,x213 }  )+$signed( { 1'b0,x214 }  )+$signed( -{ 1'b0,x215 } )+$signed( { 2'b0,x217 } <<<3'd1 )+$signed( { 2'b0,x218 } <<<3'd1 )+$signed( { 2'b0,x219 } <<<3'd1 )+$signed( -{ 1'b0,x220 } )+$signed( { 3'b0,x221 }<<<3'd2 )+$signed( -{ 2'b0,x222 }<<<3'd1 )+$signed( { 3'b0,x223 }<<<3'd2 )+$signed( -{ 2'b0,x224 }<<<3'd1 )+$signed( { 3'b0,x226 }<<<3'd2 )+$signed( -{ 2'b0,x227 }<<<3'd1 )+$signed( -{ 2'b0,x229 }<<<3'd1 )+$signed( -{ 2'b0,x230 }<<<3'd1 )+$signed( { 2'b0,x231 } <<<3'd1 )+$signed( { 2'b0,x232 } <<<3'd1 )+$signed( { 2'b0,x233 } <<<3'd1 )+$signed( -{ 1'b0,x235 } )+$signed( -{ 2'b0,x236 }<<<3'd1 )+$signed( { 3'b0,x237 }<<<3'd2 )+$signed( { 4'b0,x238 }<<<3'd3 )+$signed( -{ 2'b0,x239 }<<<3'd1 )+$signed( -{ 2'b0,x240 }<<<3'd1 )+$signed( { 1'b0,x241 }  )+$signed( { 2'b0,x243 } <<<3'd1 )+$signed( { 2'b0,x244 } <<<3'd1 )+$signed( -{ 1'b0,x245 } )+$signed( { 1'b0,x246 }  )+$signed( { 1'b0,x247 }  )+$signed( { 2'b0,x248 } <<<3'd1 )+$signed( -{ 3'b0,x249 }<<<3'd2)+$signed( -{ 1'b0,x250 } )+$signed( { 2'b0,x251 } <<<3'd1 )+$signed( -{ 3'b0,x252 }<<<3'd2)+$signed( { 1'b0,x253 }  )+$signed( { 4'b0,x255 }<<<3'd3 )+$signed( -{ 2'b0,x256 }<<<3'd1 )+$signed( -{ 3'b0,x257 }<<<3'd2)+$signed( -{ 1'b0,x260 } )+$signed( -{ 3'b0,x261 }<<<3'd2)+$signed( { 3'b0,x262 }<<<3'd2 )+$signed( { 2'b0,x265 } <<<3'd1 )+$signed( { 2'b0,x266 } <<<3'd1 )+$signed( -{ 3'b0,x268 }<<<3'd2)+$signed( -{ 2'b0,x269 }<<<3'd1 )+$signed( { 1'b0,x270 }  )+$signed( { 1'b0,x271 }  )+$signed( { 1'b0,x272 }  )+$signed( { 2'b0,x273 } <<<3'd1 )+$signed( { 1'b0,x274 }  )+$signed( -{ 2'b0,x275 }<<<3'd1 )+$signed( { 1'b0,x277 }  )+$signed( -{ 2'b0,x278 }<<<3'd1 )+$signed( -{ 1'b0,x279 } )+$signed( { 2'b0,x280 } <<<3'd1 )+$signed( -{ 1'b0,x281 } )+$signed( { 1'b0,x282 }  )+$signed( { 1'b0,x284 }  )+$signed( -{ 3'b0,x285 }<<<3'd2)+$signed( -{ 3'b0,x286 }<<<3'd2)+$signed( -{ 2'b0,x287 }<<<3'd1 )+$signed( { 2'b0,x288 } <<<3'd1 )+$signed( { 1'b0,x289 }  )+$signed( { 2'b0,x290 } <<<3'd1 )+$signed( { 3'b0,x291 }<<<3'd2 )+$signed( { 3'b0,x292 }<<<3'd2 )+$signed( { 3'b0,x293 }<<<3'd2 )+$signed( -{ 1'b0,x294 } )+$signed( { 1'b0,x295 }  )+$signed( { 2'b0,x296 } <<<3'd1 )+$signed( { 2'b0,x297 } <<<3'd1 )+$signed( -{ 1'b0,x298 } )+$signed( { 2'b0,x299 } <<<3'd1 )+$signed( -{ 3'b0,x300 }<<<3'd2)+$signed( -{ 1'b0,x301 } )+$signed( { 2'b0,x303 } <<<3'd1 )+$signed( -{ 2'b0,x304 }<<<3'd1 )+$signed( -{ 3'b0,x305 }<<<3'd2)+$signed( -{ 2'b0,x306 }<<<3'd1 )+$signed( { 3'b0,x307 }<<<3'd2 )+$signed( -{ 1'b0,x308 } )+$signed( -{ 1'b0,x309 } )+$signed( { 3'b0,x311 }<<<3'd2 )+$signed( { 2'b0,x312 } <<<3'd1 )+$signed( -{ 3'b0,x313 }<<<3'd2)+$signed( { 3'b0,x314 }<<<3'd2 )+$signed( -{ 2'b0,x315 }<<<3'd1 )+$signed( { 3'b0,x316 }<<<3'd2 )+$signed( -{ 3'b0,x318 }<<<3'd2)+$signed( -{ 1'b0,x319 } )+$signed( -{ 2'b0,x320 }<<<3'd1 )+$signed( -{ 2'b0,x321 }<<<3'd1 )+$signed( -{ 3'b0,x322 }<<<3'd2)+$signed( -{ 1'b0,x323 } )+$signed( { 3'b0,x324 }<<<3'd2 )+$signed( { 3'b0,x325 }<<<3'd2 )+$signed( { 2'b0,x327 } <<<3'd1 )+$signed( -{ 1'b0,x328 } )+$signed( -{ 1'b0,x329 } )+$signed( { 2'b0,x330 } <<<3'd1 )+$signed( -{ 4'b0, x331 }<<<3'd3 )+$signed( { 2'b0,x332 } <<<3'd1 )+$signed( { 2'b0,x333 } <<<3'd1 )+$signed( -{ 3'b0,x335 }<<<3'd2)+$signed( -{ 2'b0,x336 }<<<3'd1 )+$signed( -{ 1'b0,x339 } )+$signed( { 3'b0,x340 }<<<3'd2 )+$signed( { 2'b0,x341 } <<<3'd1 )+$signed( { 1'b0,x342 }  )+$signed( { 3'b0,x343 }<<<3'd2 )+$signed( -{ 2'b0,x344 }<<<3'd1 )+$signed( { 3'b0,x345 }<<<3'd2 )+$signed( -{ 1'b0,x346 } )+$signed( { 2'b0,x347 } <<<3'd1 )+$signed( { 1'b0,x351 }  )+$signed( -{ 1'b0,x352 } )+$signed( -{ 3'b0,x354 }<<<3'd2)+$signed( { 3'b0,x355 }<<<3'd2 )+$signed( { 1'b0,x356 }  )+$signed( -{ 1'b0,x357 } )+$signed( { 3'b0,x358 }<<<3'd2 )+$signed( { 2'b0,x360 } <<<3'd1 )+$signed( { 3'b0,x361 }<<<3'd2 )+$signed( -{ 3'b0,x362 }<<<3'd2)+$signed( -{ 1'b0,x363 } )+$signed( { 3'b0,x364 }<<<3'd2 )+$signed( { 2'b0,x365 } <<<3'd1 )+$signed( { 4'b0,x366 }<<<3'd3 )+$signed( -{ 3'b0,x367 }<<<3'd2)+$signed( { 1'b0,x368 }  )+$signed( { 1'b0,x369 }  )+$signed( { 3'b0,x370 }<<<3'd2 )+$signed( { 4'b0,x371 }<<<3'd3 )+$signed( -{ 2'b0,x372 }<<<3'd1 )+$signed( { 1'b0,x373 }  )+$signed( -{ 3'b0,x374 }<<<3'd2)+$signed( { 2'b0,x375 } <<<3'd1 )+$signed( { 2'b0,x376 } <<<3'd1 )+$signed( { 2'b0,x377 } <<<3'd1 )+$signed( { 1'b0,x378 }  )+$signed( { 3'b0,x379 }<<<3'd2 )+$signed( -{ 3'b0,x382 }<<<3'd2)+$signed( -{ 1'b0,x383 } )+$signed( { 3'b0,x384 }<<<3'd2 )+$signed( -{ 2'b0,x385 }<<<3'd1 )+$signed( -{ 1'b0,x386 } )+$signed( -{ 2'b0,x387 }<<<3'd1 )+$signed( { 2'b0,x388 } <<<3'd1 )+$signed( -{ 3'b0,x389 }<<<3'd2)+$signed( { 2'b0,x390 } <<<3'd1 )+$signed( { 2'b0,x392 } <<<3'd1 )+$signed( { 3'b0,x395 }<<<3'd2 )+$signed( { 2'b0,x396 } <<<3'd1 )+$signed( { 3'b0,x397 }<<<3'd2 )+$signed( -{ 1'b0,x398 } )+$signed( { 1'b0,x399 }  )+$signed( { 2'b0,x400 } <<<3'd1 )+$signed( -{ 2'b0,x401 }<<<3'd1 )+$signed( { 3'b0,x402 }<<<3'd2 )+$signed( -{ 2'b0,x403 }<<<3'd1 )+$signed( { 1'b0,x404 }  )+$signed( { 3'b0,x405 }<<<3'd2 )+$signed( -{ 1'b0,x406 } )+$signed( { 3'b0,x407 }<<<3'd2 )+$signed( { 4'b0,x408 }<<<3'd3 )+$signed( -{ 2'b0,x409 }<<<3'd1 )+$signed( { 2'b0,x410 } <<<3'd1 )+$signed( -{ 1'b0,x411 } )+$signed( -{ 1'b0,x412 } )+$signed( { 2'b0,x413 } <<<3'd1 )+$signed( { 2'b0,x414 } <<<3'd1 )+$signed( -{ 3'b0,x416 }<<<3'd2)+$signed( -{ 2'b0,x417 }<<<3'd1 )+$signed( { 3'b0,x418 }<<<3'd2 )+$signed( { 2'b0,x419 } <<<3'd1 )+$signed( { 3'b0,x420 }<<<3'd2 )+$signed( { 3'b0,x421 }<<<3'd2 )+$signed( { 2'b0,x423 } <<<3'd1 )+$signed( -{ 1'b0,x424 } )+$signed( -{ 2'b0,x425 }<<<3'd1 )+$signed( { 2'b0,x426 } <<<3'd1 )+$signed( { 1'b0,x427 }  )+$signed( -{ 2'b0,x428 }<<<3'd1 )+$signed( -{ 1'b0,x429 } )+$signed( { 3'b0,x430 }<<<3'd2 )+$signed( { 2'b0,x431 } <<<3'd1 )+$signed( { 1'b0,x432 }  )+$signed( -{ 2'b0,x433 }<<<3'd1 )+$signed( -{ 1'b0,x434 } )+$signed( -{ 1'b0,x436 } )+$signed( -{ 1'b0,x437 } )+$signed( -{ 1'b0,x438 } )+$signed( { 3'b0,x439 }<<<3'd2 )+$signed( -{ 2'b0,x440 }<<<3'd1 )+$signed( -{ 2'b0,x441 }<<<3'd1 )+$signed( { 3'b0,x443 }<<<3'd2 )+$signed( { 3'b0,x444 }<<<3'd2 )+$signed( -{ 2'b0,x445 }<<<3'd1 )+$signed( { 2'b0,x446 } <<<3'd1 )+$signed( -{ 2'b0,x449 }<<<3'd1 )+$signed( -{ 2'b0,x450 }<<<3'd1 )+$signed( -{ 1'b0,x451 } )+$signed( -{ 3'b0,x452 }<<<3'd2)+$signed( -{ 1'b0,x453 } )+$signed( -{ 3'b0,x454 }<<<3'd2)+$signed( -{ 1'b0,x455 } )+$signed( { 2'b0,x456 } <<<3'd1 )+$signed( { 3'b0,x457 }<<<3'd2 )+$signed( -{ 2'b0,x458 }<<<3'd1 )+$signed( { 2'b0,x459 } <<<3'd1 )+$signed( { 2'b0,x460 } <<<3'd1 )+$signed( { 1'b0,x462 }  )+$signed( -{ 2'b0,x463 }<<<3'd1 )+$signed( -{ 3'b0,x464 }<<<3'd2)+$signed( -{ 3'b0,x465 }<<<3'd2)+$signed( { 2'b0,x466 } <<<3'd1 )+$signed( -{ 2'b0,x467 }<<<3'd1 )+$signed( { 3'b0,x468 }<<<3'd2 )+$signed( -{ 1'b0,x469 } )+$signed( { 3'b0,x470 }<<<3'd2 )+$signed( -{ 3'b0,x471 }<<<3'd2)+$signed( { 2'b0,x472 } <<<3'd1 )+$signed( -{ 3'b0,x474 }<<<3'd2)+$signed( { 1'b0,x475 }  )+$signed( -{ 2'b0,x476 }<<<3'd1 )+$signed( -{ 2'b0,x477 }<<<3'd1 )+$signed( -{ 3'b0,x478 }<<<3'd2)+$signed( { 2'b0,x479 } <<<3'd1 )+$signed( { 3'b0,x481 }<<<3'd2 )+$signed( { 2'b0,x482 } <<<3'd1 )+$signed( { 3'b0,x483 }<<<3'd2 )+$signed( { 2'b0,x485 } <<<3'd1 )+$signed( -{ 2'b0,x486 }<<<3'd1 )+$signed( -{ 2'b0,x487 }<<<3'd1 )+$signed( -{ 3'b0,x488 }<<<3'd2)+$signed( -{ 2'b0,x489 }<<<3'd1 )+$signed( -{ 2'b0,x490 }<<<3'd1 )+$signed( { 1'b0,x491 }  )+$signed( -{ 2'b0,x492 }<<<3'd1 )+$signed( -{ 3'b0,x493 }<<<3'd2)+$signed( { 1'b0,x494 }  )-$signed(13'd8);
assign y13=temp_y[13][13] ==1'b1 ? 6'd0 :  
    temp_y[13][10] ==1'b1 ? 6'd63 : 
    temp_y[13][3]==1'b1 ? temp_y[13][9:4]+1'b1 : temp_y[13][9:4];
assign temp_y[14] = 
+$signed( { 2'b0,x2 } <<<3'd1 )+$signed( { 2'b0,x3 } <<<3'd1 )+$signed( -{ 2'b0,x4 }<<<3'd1 )+$signed( { 1'b0,x5 }  )+$signed( { 1'b0,x6 }  )+$signed( -{ 2'b0,x7 }<<<3'd1 )+$signed( -{ 3'b0,x8 }<<<3'd2)+$signed( { 2'b0,x9 } <<<3'd1 )+$signed( { 2'b0,x10 } <<<3'd1 )+$signed( { 2'b0,x11 } <<<3'd1 )+$signed( -{ 1'b0,x14 } )+$signed( -{ 3'b0,x15 }<<<3'd2)+$signed( { 1'b0,x16 }  )+$signed( { 1'b0,x19 }  )+$signed( -{ 3'b0,x20 }<<<3'd2)+$signed( { 3'b0,x21 }<<<3'd2 )+$signed( -{ 1'b0,x22 } )+$signed( { 3'b0,x23 }<<<3'd2 )+$signed( { 2'b0,x24 } <<<3'd1 )+$signed( { 1'b0,x25 }  )+$signed( -{ 3'b0,x26 }<<<3'd2)+$signed( { 2'b0,x28 } <<<3'd1 )+$signed( -{ 1'b0,x29 } )+$signed( -{ 3'b0,x30 }<<<3'd2)+$signed( { 1'b0,x31 }  )+$signed( { 3'b0,x32 }<<<3'd2 )+$signed( -{ 3'b0,x33 }<<<3'd2)+$signed( { 2'b0,x34 } <<<3'd1 )+$signed( { 1'b0,x35 }  )+$signed( -{ 3'b0,x36 }<<<3'd2)+$signed( -{ 2'b0,x37 }<<<3'd1 )+$signed( -{ 2'b0,x38 }<<<3'd1 )+$signed( { 3'b0,x39 }<<<3'd2 )+$signed( { 1'b0,x40 }  )+$signed( { 1'b0,x41 }  )+$signed( -{ 2'b0,x42 }<<<3'd1 )+$signed( { 2'b0,x43 } <<<3'd1 )+$signed( -{ 2'b0,x44 }<<<3'd1 )+$signed( { 1'b0,x45 }  )+$signed( { 1'b0,x46 }  )+$signed( -{ 2'b0,x47 }<<<3'd1 )+$signed( { 1'b0,x48 }  )+$signed( -{ 1'b0,x49 } )+$signed( { 2'b0,x50 } <<<3'd1 )+$signed( { 2'b0,x52 } <<<3'd1 )+$signed( -{ 2'b0,x53 }<<<3'd1 )+$signed( -{ 2'b0,x54 }<<<3'd1 )+$signed( -{ 2'b0,x55 }<<<3'd1 )+$signed( -{ 1'b0,x56 } )+$signed( { 3'b0,x57 }<<<3'd2 )+$signed( { 1'b0,x58 }  )+$signed( -{ 1'b0,x59 } )+$signed( -{ 2'b0,x60 }<<<3'd1 )+$signed( -{ 1'b0,x61 } )+$signed( -{ 3'b0,x62 }<<<3'd2)+$signed( { 2'b0,x64 } <<<3'd1 )+$signed( { 1'b0,x66 }  )+$signed( -{ 2'b0,x67 }<<<3'd1 )+$signed( -{ 3'b0,x68 }<<<3'd2)+$signed( -{ 3'b0,x69 }<<<3'd2)+$signed( { 3'b0,x70 }<<<3'd2 )+$signed( { 1'b0,x71 }  )+$signed( -{ 3'b0,x72 }<<<3'd2)+$signed( { 1'b0,x73 }  )+$signed( { 2'b0,x74 } <<<3'd1 )+$signed( { 3'b0,x75 }<<<3'd2 )+$signed( -{ 2'b0,x76 }<<<3'd1 )+$signed( { 1'b0,x77 }  )+$signed( { 3'b0,x78 }<<<3'd2 )+$signed( { 2'b0,x79 } <<<3'd1 )+$signed( { 1'b0,x80 }  )+$signed( -{ 1'b0,x81 } )+$signed( -{ 1'b0,x82 } )+$signed( -{ 3'b0,x84 }<<<3'd2)+$signed( -{ 2'b0,x85 }<<<3'd1 )+$signed( -{ 3'b0,x86 }<<<3'd2)+$signed( { 1'b0,x87 }  )+$signed( -{ 1'b0,x91 } )+$signed( { 4'b0,x93 }<<<3'd3 )+$signed( -{ 1'b0,x94 } )+$signed( { 1'b0,x96 }  )+$signed( { 2'b0,x98 } <<<3'd1 )+$signed( -{ 4'b0, x99 }<<<3'd3 )+$signed( -{ 1'b0,x100 } )+$signed( -{ 2'b0,x101 }<<<3'd1 )+$signed( { 2'b0,x102 } <<<3'd1 )+$signed( -{ 2'b0,x103 }<<<3'd1 )+$signed( { 2'b0,x104 } <<<3'd1 )+$signed( -{ 1'b0,x105 } )+$signed( -{ 3'b0,x107 }<<<3'd2)+$signed( -{ 3'b0,x108 }<<<3'd2)+$signed( -{ 2'b0,x109 }<<<3'd1 )+$signed( { 2'b0,x110 } <<<3'd1 )+$signed( { 3'b0,x111 }<<<3'd2 )+$signed( -{ 1'b0,x112 } )+$signed( -{ 3'b0,x113 }<<<3'd2)+$signed( { 2'b0,x114 } <<<3'd1 )+$signed( { 3'b0,x115 }<<<3'd2 )+$signed( { 2'b0,x116 } <<<3'd1 )+$signed( -{ 3'b0,x117 }<<<3'd2)+$signed( -{ 1'b0,x118 } )+$signed( -{ 2'b0,x119 }<<<3'd1 )+$signed( { 2'b0,x120 } <<<3'd1 )+$signed( -{ 2'b0,x121 }<<<3'd1 )+$signed( { 1'b0,x123 }  )+$signed( -{ 3'b0,x124 }<<<3'd2)+$signed( -{ 2'b0,x125 }<<<3'd1 )+$signed( { 1'b0,x127 }  )+$signed( -{ 2'b0,x128 }<<<3'd1 )+$signed( { 1'b0,x129 }  )+$signed( -{ 2'b0,x130 }<<<3'd1 )+$signed( { 2'b0,x131 } <<<3'd1 )+$signed( { 2'b0,x132 } <<<3'd1 )+$signed( { 3'b0,x133 }<<<3'd2 )+$signed( -{ 3'b0,x135 }<<<3'd2)+$signed( -{ 1'b0,x136 } )+$signed( { 2'b0,x137 } <<<3'd1 )+$signed( -{ 2'b0,x140 }<<<3'd1 )+$signed( { 1'b0,x141 }  )+$signed( { 2'b0,x142 } <<<3'd1 )+$signed( { 3'b0,x143 }<<<3'd2 )+$signed( { 3'b0,x144 }<<<3'd2 )+$signed( { 2'b0,x145 } <<<3'd1 )+$signed( -{ 2'b0,x146 }<<<3'd1 )+$signed( -{ 4'b0, x147 }<<<3'd3 )+$signed( -{ 3'b0,x148 }<<<3'd2)+$signed( -{ 2'b0,x149 }<<<3'd1 )+$signed( -{ 3'b0,x151 }<<<3'd2)+$signed( -{ 3'b0,x152 }<<<3'd2)+$signed( { 1'b0,x153 }  )+$signed( { 2'b0,x156 } <<<3'd1 )+$signed( { 1'b0,x157 }  )+$signed( -{ 3'b0,x158 }<<<3'd2)+$signed( { 3'b0,x159 }<<<3'd2 )+$signed( -{ 3'b0,x160 }<<<3'd2)+$signed( { 2'b0,x161 } <<<3'd1 )+$signed( { 2'b0,x162 } <<<3'd1 )+$signed( { 2'b0,x164 } <<<3'd1 )+$signed( -{ 4'b0, x165 }<<<3'd3 )+$signed( -{ 2'b0,x167 }<<<3'd1 )+$signed( { 1'b0,x168 }  )+$signed( -{ 4'b0, x169 }<<<3'd3 )+$signed( { 4'b0,x170 }<<<3'd3 )+$signed( { 2'b0,x172 } <<<3'd1 )+$signed( { 3'b0,x173 }<<<3'd2 )+$signed( -{ 3'b0,x174 }<<<3'd2)+$signed( -{ 1'b0,x175 } )+$signed( -{ 2'b0,x177 }<<<3'd1 )+$signed( -{ 2'b0,x178 }<<<3'd1 )+$signed( { 3'b0,x179 }<<<3'd2 )+$signed( -{ 2'b0,x180 }<<<3'd1 )+$signed( { 2'b0,x182 } <<<3'd1 )+$signed( -{ 4'b0, x183 }<<<3'd3 )+$signed( -{ 3'b0,x184 }<<<3'd2)+$signed( { 3'b0,x186 }<<<3'd2 )+$signed( -{ 4'b0, x187 }<<<3'd3 )+$signed( { 4'b0,x188 }<<<3'd3 )+$signed( { 2'b0,x189 } <<<3'd1 )+$signed( { 3'b0,x190 }<<<3'd2 )+$signed( { 3'b0,x191 }<<<3'd2 )+$signed( -{ 3'b0,x192 }<<<3'd2)+$signed( -{ 1'b0,x193 } )+$signed( -{ 2'b0,x194 }<<<3'd1 )+$signed( { 1'b0,x195 }  )+$signed( -{ 1'b0,x196 } )+$signed( { 3'b0,x197 }<<<3'd2 )+$signed( -{ 2'b0,x198 }<<<3'd1 )+$signed( -{ 3'b0,x200 }<<<3'd2)+$signed( { 1'b0,x201 }  )+$signed( -{ 2'b0,x202 }<<<3'd1 )+$signed( { 2'b0,x203 } <<<3'd1 )+$signed( { 3'b0,x204 }<<<3'd2 )+$signed( -{ 4'b0, x205 }<<<3'd3 )+$signed( { 1'b0,x206 }  )+$signed( -{ 1'b0,x207 } )+$signed( { 2'b0,x208 } <<<3'd1 )+$signed( -{ 1'b0,x209 } )+$signed( { 3'b0,x210 }<<<3'd2 )+$signed( -{ 2'b0,x212 }<<<3'd1 )+$signed( { 2'b0,x214 } <<<3'd1 )+$signed( { 3'b0,x215 }<<<3'd2 )+$signed( { 1'b0,x216 }  )+$signed( -{ 3'b0,x217 }<<<3'd2)+$signed( { 4'b0,x218 }<<<3'd3 )+$signed( -{ 1'b0,x219 } )+$signed( -{ 2'b0,x220 }<<<3'd1 )+$signed( -{ 2'b0,x221 }<<<3'd1 )+$signed( -{ 2'b0,x222 }<<<3'd1 )+$signed( -{ 3'b0,x224 }<<<3'd2)+$signed( -{ 1'b0,x225 } )+$signed( { 1'b0,x226 }  )+$signed( { 2'b0,x227 } <<<3'd1 )+$signed( { 2'b0,x228 } <<<3'd1 )+$signed( -{ 1'b0,x229 } )+$signed( { 2'b0,x230 } <<<3'd1 )+$signed( -{ 2'b0,x231 }<<<3'd1 )+$signed( { 4'b0,x232 }<<<3'd3 )+$signed( -{ 3'b0,x233 }<<<3'd2)+$signed( -{ 1'b0,x234 } )+$signed( -{ 2'b0,x235 }<<<3'd1 )+$signed( { 4'b0,x236 }<<<3'd3 )+$signed( -{ 3'b0,x237 }<<<3'd2)+$signed( { 1'b0,x238 }  )+$signed( -{ 3'b0,x239 }<<<3'd2)+$signed( -{ 1'b0,x240 } )+$signed( -{ 3'b0,x242 }<<<3'd2)+$signed( { 2'b0,x243 } <<<3'd1 )+$signed( -{ 3'b0,x244 }<<<3'd2)+$signed( { 1'b0,x245 }  )+$signed( { 3'b0,x246 }<<<3'd2 )+$signed( { 2'b0,x247 } <<<3'd1 )+$signed( -{ 2'b0,x248 }<<<3'd1 )+$signed( { 3'b0,x249 }<<<3'd2 )+$signed( { 1'b0,x250 }  )+$signed( -{ 4'b0, x251 }<<<3'd3 )+$signed( { 2'b0,x254 } <<<3'd1 )+$signed( -{ 3'b0,x255 }<<<3'd2)+$signed( { 2'b0,x256 } <<<3'd1 )+$signed( -{ 3'b0,x257 }<<<3'd2)+$signed( -{ 1'b0,x258 } )+$signed( -{ 1'b0,x259 } )+$signed( -{ 2'b0,x260 }<<<3'd1 )+$signed( { 3'b0,x261 }<<<3'd2 )+$signed( -{ 4'b0, x262 }<<<3'd3 )+$signed( { 2'b0,x263 } <<<3'd1 )+$signed( { 3'b0,x264 }<<<3'd2 )+$signed( { 2'b0,x265 } <<<3'd1 )+$signed( -{ 2'b0,x266 }<<<3'd1 )+$signed( { 1'b0,x267 }  )+$signed( { 3'b0,x268 }<<<3'd2 )+$signed( -{ 1'b0,x269 } )+$signed( { 2'b0,x270 } <<<3'd1 )+$signed( -{ 1'b0,x271 } )+$signed( { 3'b0,x272 }<<<3'd2 )+$signed( -{ 4'b0, x273 }<<<3'd3 )+$signed( { 1'b0,x274 }  )+$signed( -{ 2'b0,x275 }<<<3'd1 )+$signed( -{ 2'b0,x276 }<<<3'd1 )+$signed( { 4'b0,x277 }<<<3'd3 )+$signed( -{ 3'b0,x278 }<<<3'd2)+$signed( { 1'b0,x279 }  )+$signed( { 3'b0,x281 }<<<3'd2 )+$signed( { 1'b0,x282 }  )+$signed( { 1'b0,x284 }  )+$signed( { 3'b0,x285 }<<<3'd2 )+$signed( { 2'b0,x286 } <<<3'd1 )+$signed( -{ 3'b0,x287 }<<<3'd2)+$signed( -{ 3'b0,x288 }<<<3'd2)+$signed( -{ 2'b0,x289 }<<<3'd1 )+$signed( { 3'b0,x290 }<<<3'd2 )+$signed( -{ 3'b0,x291 }<<<3'd2)+$signed( { 2'b0,x292 } <<<3'd1 )+$signed( -{ 3'b0,x293 }<<<3'd2)+$signed( -{ 1'b0,x294 } )+$signed( -{ 3'b0,x295 }<<<3'd2)+$signed( { 1'b0,x296 }  )+$signed( -{ 3'b0,x297 }<<<3'd2)+$signed( -{ 3'b0,x298 }<<<3'd2)+$signed( -{ 3'b0,x299 }<<<3'd2)+$signed( { 2'b0,x301 } <<<3'd1 )+$signed( -{ 2'b0,x302 }<<<3'd1 )+$signed( { 1'b0,x303 }  )+$signed( { 3'b0,x304 }<<<3'd2 )+$signed( -{ 3'b0,x305 }<<<3'd2)+$signed( { 3'b0,x309 }<<<3'd2 )+$signed( -{ 1'b0,x310 } )+$signed( { 1'b0,x311 }  )+$signed( -{ 2'b0,x312 }<<<3'd1 )+$signed( { 3'b0,x313 }<<<3'd2 )+$signed( { 2'b0,x314 } <<<3'd1 )+$signed( -{ 2'b0,x315 }<<<3'd1 )+$signed( { 3'b0,x316 }<<<3'd2 )+$signed( -{ 3'b0,x317 }<<<3'd2)+$signed( -{ 1'b0,x318 } )+$signed( -{ 3'b0,x319 }<<<3'd2)+$signed( -{ 1'b0,x320 } )+$signed( -{ 3'b0,x321 }<<<3'd2)+$signed( -{ 1'b0,x322 } )+$signed( -{ 3'b0,x323 }<<<3'd2)+$signed( -{ 3'b0,x324 }<<<3'd2)+$signed( { 3'b0,x327 }<<<3'd2 )+$signed( -{ 2'b0,x328 }<<<3'd1 )+$signed( { 2'b0,x329 } <<<3'd1 )+$signed( -{ 3'b0,x330 }<<<3'd2)+$signed( -{ 1'b0,x331 } )+$signed( -{ 1'b0,x332 } )+$signed( -{ 2'b0,x333 }<<<3'd1 )+$signed( { 1'b0,x334 }  )+$signed( { 1'b0,x336 }  )+$signed( -{ 2'b0,x338 }<<<3'd1 )+$signed( -{ 1'b0,x339 } )+$signed( -{ 3'b0,x340 }<<<3'd2)+$signed( -{ 1'b0,x341 } )+$signed( { 2'b0,x342 } <<<3'd1 )+$signed( -{ 2'b0,x343 }<<<3'd1 )+$signed( -{ 3'b0,x344 }<<<3'd2)+$signed( { 2'b0,x345 } <<<3'd1 )+$signed( { 2'b0,x346 } <<<3'd1 )+$signed( { 3'b0,x348 }<<<3'd2 )+$signed( { 3'b0,x349 }<<<3'd2 )+$signed( -{ 2'b0,x350 }<<<3'd1 )+$signed( -{ 1'b0,x351 } )+$signed( { 2'b0,x354 } <<<3'd1 )+$signed( { 3'b0,x355 }<<<3'd2 )+$signed( { 1'b0,x356 }  )+$signed( { 1'b0,x357 }  )+$signed( { 2'b0,x358 } <<<3'd1 )+$signed( { 1'b0,x359 }  )+$signed( -{ 2'b0,x360 }<<<3'd1 )+$signed( -{ 1'b0,x361 } )+$signed( { 3'b0,x362 }<<<3'd2 )+$signed( { 1'b0,x363 }  )+$signed( { 4'b0,x364 }<<<3'd3 )+$signed( -{ 1'b0,x365 } )+$signed( -{ 1'b0,x366 } )+$signed( -{ 2'b0,x369 }<<<3'd1 )+$signed( { 2'b0,x370 } <<<3'd1 )+$signed( { 3'b0,x371 }<<<3'd2 )+$signed( { 1'b0,x372 }  )+$signed( -{ 2'b0,x373 }<<<3'd1 )+$signed( -{ 2'b0,x374 }<<<3'd1 )+$signed( { 3'b0,x375 }<<<3'd2 )+$signed( -{ 2'b0,x376 }<<<3'd1 )+$signed( { 4'b0,x377 }<<<3'd3 )+$signed( { 1'b0,x378 }  )+$signed( -{ 3'b0,x379 }<<<3'd2)+$signed( -{ 3'b0,x380 }<<<3'd2)+$signed( { 1'b0,x381 }  )+$signed( -{ 2'b0,x382 }<<<3'd1 )+$signed( -{ 3'b0,x383 }<<<3'd2)+$signed( { 1'b0,x384 }  )+$signed( -{ 2'b0,x385 }<<<3'd1 )+$signed( -{ 2'b0,x386 }<<<3'd1 )+$signed( -{ 1'b0,x387 } )+$signed( -{ 2'b0,x388 }<<<3'd1 )+$signed( { 3'b0,x389 }<<<3'd2 )+$signed( { 2'b0,x390 } <<<3'd1 )+$signed( { 3'b0,x391 }<<<3'd2 )+$signed( { 3'b0,x392 }<<<3'd2 )+$signed( -{ 2'b0,x393 }<<<3'd1 )+$signed( -{ 1'b0,x394 } )+$signed( -{ 2'b0,x395 }<<<3'd1 )+$signed( -{ 3'b0,x396 }<<<3'd2)+$signed( -{ 2'b0,x397 }<<<3'd1 )+$signed( -{ 3'b0,x398 }<<<3'd2)+$signed( -{ 3'b0,x399 }<<<3'd2)+$signed( { 3'b0,x401 }<<<3'd2 )+$signed( { 1'b0,x402 }  )+$signed( -{ 4'b0, x403 }<<<3'd3 )+$signed( -{ 3'b0,x404 }<<<3'd2)+$signed( -{ 1'b0,x405 } )+$signed( { 1'b0,x406 }  )+$signed( { 3'b0,x407 }<<<3'd2 )+$signed( { 3'b0,x408 }<<<3'd2 )+$signed( -{ 3'b0,x409 }<<<3'd2)+$signed( -{ 1'b0,x410 } )+$signed( { 2'b0,x412 } <<<3'd1 )+$signed( -{ 3'b0,x413 }<<<3'd2)+$signed( { 4'b0,x414 }<<<3'd3 )+$signed( { 3'b0,x415 }<<<3'd2 )+$signed( -{ 4'b0, x416 }<<<3'd3 )+$signed( -{ 3'b0,x417 }<<<3'd2)+$signed( -{ 2'b0,x418 }<<<3'd1 )+$signed( -{ 2'b0,x419 }<<<3'd1 )+$signed( -{ 1'b0,x420 } )+$signed( { 2'b0,x421 } <<<3'd1 )+$signed( { 3'b0,x422 }<<<3'd2 )+$signed( { 2'b0,x423 } <<<3'd1 )+$signed( { 3'b0,x424 }<<<3'd2 )+$signed( { 1'b0,x425 }  )+$signed( -{ 3'b0,x426 }<<<3'd2)+$signed( { 3'b0,x427 }<<<3'd2 )+$signed( -{ 1'b0,x428 } )+$signed( { 4'b0,x429 }<<<3'd3 )+$signed( -{ 3'b0,x430 }<<<3'd2)+$signed( -{ 3'b0,x431 }<<<3'd2)+$signed( { 3'b0,x432 }<<<3'd2 )+$signed( { 3'b0,x433 }<<<3'd2 )+$signed( { 4'b0,x434 }<<<3'd3 )+$signed( { 4'b0,x435 }<<<3'd3 )+$signed( { 2'b0,x436 } <<<3'd1 )+$signed( { 1'b0,x437 }  )+$signed( -{ 4'b0, x439 }<<<3'd3 )+$signed( -{ 1'b0,x440 } )+$signed( -{ 2'b0,x441 }<<<3'd1 )+$signed( -{ 3'b0,x442 }<<<3'd2)+$signed( -{ 3'b0,x443 }<<<3'd2)+$signed( -{ 1'b0,x444 } )+$signed( { 4'b0,x445 }<<<3'd3 )+$signed( -{ 3'b0,x446 }<<<3'd2)+$signed( { 3'b0,x447 }<<<3'd2 )+$signed( -{ 3'b0,x448 }<<<3'd2)+$signed( { 3'b0,x449 }<<<3'd2 )+$signed( { 2'b0,x450 } <<<3'd1 )+$signed( { 2'b0,x451 } <<<3'd1 )+$signed( { 4'b0,x452 }<<<3'd3 )+$signed( -{ 1'b0,x453 } )+$signed( { 3'b0,x454 }<<<3'd2 )+$signed( -{ 5'b0,x455 }<<<3'd4 )+$signed( -{ 3'b0,x457 }<<<3'd2)+$signed( { 2'b0,x459 } <<<3'd1 )+$signed( { 1'b0,x460 }  )+$signed( -{ 3'b0,x461 }<<<3'd2)+$signed( { 3'b0,x462 }<<<3'd2 )+$signed( { 4'b0,x463 }<<<3'd3 )+$signed( { 2'b0,x464 } <<<3'd1 )+$signed( { 4'b0,x465 }<<<3'd3 )+$signed( -{ 1'b0,x466 } )+$signed( { 4'b0,x467 }<<<3'd3 )+$signed( -{ 1'b0,x468 } )+$signed( -{ 4'b0, x469 }<<<3'd3 )+$signed( -{ 2'b0,x470 }<<<3'd1 )+$signed( -{ 4'b0, x472 }<<<3'd3 )+$signed( { 1'b0,x473 }  )+$signed( -{ 3'b0,x474 }<<<3'd2)+$signed( { 2'b0,x475 } <<<3'd1 )+$signed( { 4'b0,x476 }<<<3'd3 )+$signed( { 1'b0,x477 }  )+$signed( { 4'b0,x478 }<<<3'd3 )+$signed( -{ 1'b0,x479 } )+$signed( { 4'b0,x480 }<<<3'd3 )+$signed( -{ 3'b0,x481 }<<<3'd2)+$signed( { 3'b0,x482 }<<<3'd2 )+$signed( { 2'b0,x483 } <<<3'd1 )+$signed( -{ 2'b0,x484 }<<<3'd1 )+$signed( -{ 4'b0, x485 }<<<3'd3 )+$signed( { 4'b0,x486 }<<<3'd3 )+$signed( { 2'b0,x487 } <<<3'd1 )+$signed( { 3'b0,x488 }<<<3'd2 )+$signed( { 3'b0,x489 }<<<3'd2 )+$signed( { 4'b0,x490 }<<<3'd3 )+$signed( { 2'b0,x491 } <<<3'd1 )+$signed( { 2'b0,x492 } <<<3'd1 )+$signed( { 3'b0,x493 }<<<3'd2 )+$signed( -{ 3'b0,x494 }<<<3'd2)+$signed( { 3'b0,x495 }<<<3'd2 )-$signed(13'd8);
assign y14=temp_y[14][13] ==1'b1 ? 6'd0 :  
    temp_y[14][10] ==1'b1 ? 6'd63 : 
    temp_y[14][3]==1'b1 ? temp_y[14][9:4]+1'b1 : temp_y[14][9:4];
assign temp_y[15] = 
+$signed( -{ 3'b0,x0 }<<<3'd2)+$signed( -{ 2'b0,x1 }<<<3'd1 )+$signed( { 2'b0,x2 } <<<3'd1 )+$signed( { 2'b0,x3 } <<<3'd1 )+$signed( { 1'b0,x4 }  )+$signed( { 1'b0,x6 }  )+$signed( -{ 1'b0,x7 } )+$signed( -{ 4'b0, x8 }<<<3'd3 )+$signed( -{ 2'b0,x9 }<<<3'd1 )+$signed( { 3'b0,x10 }<<<3'd2 )+$signed( -{ 1'b0,x11 } )+$signed( -{ 3'b0,x12 }<<<3'd2)+$signed( -{ 2'b0,x13 }<<<3'd1 )+$signed( { 2'b0,x14 } <<<3'd1 )+$signed( { 1'b0,x15 }  )+$signed( { 2'b0,x16 } <<<3'd1 )+$signed( -{ 1'b0,x17 } )+$signed( -{ 3'b0,x18 }<<<3'd2)+$signed( -{ 3'b0,x19 }<<<3'd2)+$signed( -{ 3'b0,x20 }<<<3'd2)+$signed( { 2'b0,x21 } <<<3'd1 )+$signed( { 2'b0,x22 } <<<3'd1 )+$signed( { 3'b0,x23 }<<<3'd2 )+$signed( { 2'b0,x24 } <<<3'd1 )+$signed( -{ 1'b0,x25 } )+$signed( -{ 3'b0,x26 }<<<3'd2)+$signed( -{ 1'b0,x27 } )+$signed( { 3'b0,x28 }<<<3'd2 )+$signed( -{ 4'b0, x30 }<<<3'd3 )+$signed( { 1'b0,x31 }  )+$signed( -{ 3'b0,x32 }<<<3'd2)+$signed( { 1'b0,x33 }  )+$signed( -{ 3'b0,x34 }<<<3'd2)+$signed( -{ 2'b0,x36 }<<<3'd1 )+$signed( -{ 2'b0,x37 }<<<3'd1 )+$signed( { 2'b0,x38 } <<<3'd1 )+$signed( { 3'b0,x39 }<<<3'd2 )+$signed( { 2'b0,x40 } <<<3'd1 )+$signed( { 2'b0,x41 } <<<3'd1 )+$signed( { 3'b0,x42 }<<<3'd2 )+$signed( { 3'b0,x43 }<<<3'd2 )+$signed( -{ 4'b0, x44 }<<<3'd3 )+$signed( -{ 3'b0,x45 }<<<3'd2)+$signed( { 3'b0,x46 }<<<3'd2 )+$signed( -{ 4'b0, x48 }<<<3'd3 )+$signed( -{ 2'b0,x49 }<<<3'd1 )+$signed( -{ 1'b0,x50 } )+$signed( -{ 3'b0,x51 }<<<3'd2)+$signed( { 2'b0,x52 } <<<3'd1 )+$signed( -{ 2'b0,x53 }<<<3'd1 )+$signed( -{ 1'b0,x55 } )+$signed( { 1'b0,x56 }  )+$signed( { 1'b0,x57 }  )+$signed( { 1'b0,x58 }  )+$signed( -{ 2'b0,x59 }<<<3'd1 )+$signed( -{ 1'b0,x60 } )+$signed( -{ 2'b0,x61 }<<<3'd1 )+$signed( -{ 4'b0, x62 }<<<3'd3 )+$signed( -{ 2'b0,x63 }<<<3'd1 )+$signed( { 3'b0,x64 }<<<3'd2 )+$signed( -{ 3'b0,x66 }<<<3'd2)+$signed( -{ 2'b0,x67 }<<<3'd1 )+$signed( { 3'b0,x70 }<<<3'd2 )+$signed( -{ 2'b0,x71 }<<<3'd1 )+$signed( -{ 3'b0,x72 }<<<3'd2)+$signed( -{ 3'b0,x73 }<<<3'd2)+$signed( { 1'b0,x74 }  )+$signed( { 1'b0,x75 }  )+$signed( -{ 3'b0,x76 }<<<3'd2)+$signed( { 2'b0,x78 } <<<3'd1 )+$signed( { 3'b0,x79 }<<<3'd2 )+$signed( -{ 4'b0, x80 }<<<3'd3 )+$signed( { 2'b0,x81 } <<<3'd1 )+$signed( -{ 1'b0,x83 } )+$signed( { 3'b0,x84 }<<<3'd2 )+$signed( { 1'b0,x85 }  )+$signed( { 2'b0,x86 } <<<3'd1 )+$signed( { 2'b0,x87 } <<<3'd1 )+$signed( { 1'b0,x88 }  )+$signed( -{ 2'b0,x91 }<<<3'd1 )+$signed( -{ 3'b0,x92 }<<<3'd2)+$signed( { 3'b0,x93 }<<<3'd2 )+$signed( -{ 2'b0,x94 }<<<3'd1 )+$signed( -{ 4'b0, x95 }<<<3'd3 )+$signed( { 2'b0,x96 } <<<3'd1 )+$signed( { 3'b0,x97 }<<<3'd2 )+$signed( { 3'b0,x98 }<<<3'd2 )+$signed( -{ 3'b0,x99 }<<<3'd2)+$signed( { 2'b0,x100 } <<<3'd1 )+$signed( { 1'b0,x102 }  )+$signed( { 2'b0,x103 } <<<3'd1 )+$signed( -{ 2'b0,x104 }<<<3'd1 )+$signed( { 2'b0,x105 } <<<3'd1 )+$signed( -{ 1'b0,x106 } )+$signed( { 1'b0,x107 }  )+$signed( { 3'b0,x108 }<<<3'd2 )+$signed( -{ 1'b0,x109 } )+$signed( { 1'b0,x110 }  )+$signed( { 4'b0,x111 }<<<3'd3 )+$signed( -{ 3'b0,x112 }<<<3'd2)+$signed( -{ 4'b0, x113 }<<<3'd3 )+$signed( { 3'b0,x114 }<<<3'd2 )+$signed( { 3'b0,x115 }<<<3'd2 )+$signed( { 4'b0,x116 }<<<3'd3 )+$signed( -{ 4'b0, x117 }<<<3'd3 )+$signed( { 3'b0,x118 }<<<3'd2 )+$signed( -{ 3'b0,x119 }<<<3'd2)+$signed( { 3'b0,x120 }<<<3'd2 )+$signed( { 1'b0,x121 }  )+$signed( -{ 2'b0,x122 }<<<3'd1 )+$signed( -{ 2'b0,x123 }<<<3'd1 )+$signed( { 3'b0,x124 }<<<3'd2 )+$signed( { 3'b0,x125 }<<<3'd2 )+$signed( { 3'b0,x126 }<<<3'd2 )+$signed( { 1'b0,x127 }  )+$signed( { 3'b0,x128 }<<<3'd2 )+$signed( -{ 1'b0,x130 } )+$signed( -{ 1'b0,x131 } )+$signed( -{ 1'b0,x132 } )+$signed( -{ 1'b0,x133 } )+$signed( -{ 4'b0, x134 }<<<3'd3 )+$signed( { 1'b0,x135 }  )+$signed( -{ 1'b0,x136 } )+$signed( { 2'b0,x139 } <<<3'd1 )+$signed( -{ 2'b0,x140 }<<<3'd1 )+$signed( { 3'b0,x141 }<<<3'd2 )+$signed( { 3'b0,x142 }<<<3'd2 )+$signed( -{ 3'b0,x143 }<<<3'd2)+$signed( { 2'b0,x145 } <<<3'd1 )+$signed( -{ 2'b0,x146 }<<<3'd1 )+$signed( { 2'b0,x147 } <<<3'd1 )+$signed( -{ 3'b0,x148 }<<<3'd2)+$signed( { 4'b0,x149 }<<<3'd3 )+$signed( -{ 2'b0,x151 }<<<3'd1 )+$signed( -{ 2'b0,x152 }<<<3'd1 )+$signed( -{ 3'b0,x153 }<<<3'd2)+$signed( { 2'b0,x154 } <<<3'd1 )+$signed( { 1'b0,x155 }  )+$signed( { 3'b0,x156 }<<<3'd2 )+$signed( { 1'b0,x157 }  )+$signed( { 3'b0,x158 }<<<3'd2 )+$signed( { 2'b0,x159 } <<<3'd1 )+$signed( -{ 2'b0,x160 }<<<3'd1 )+$signed( { 3'b0,x161 }<<<3'd2 )+$signed( -{ 3'b0,x162 }<<<3'd2)+$signed( -{ 2'b0,x163 }<<<3'd1 )+$signed( { 1'b0,x164 }  )+$signed( -{ 1'b0,x165 } )+$signed( -{ 1'b0,x166 } )+$signed( -{ 1'b0,x167 } )+$signed( { 1'b0,x168 }  )+$signed( { 1'b0,x169 }  )+$signed( { 3'b0,x170 }<<<3'd2 )+$signed( -{ 3'b0,x171 }<<<3'd2)+$signed( -{ 3'b0,x172 }<<<3'd2)+$signed( -{ 1'b0,x173 } )+$signed( -{ 2'b0,x174 }<<<3'd1 )+$signed( -{ 1'b0,x175 } )+$signed( { 2'b0,x176 } <<<3'd1 )+$signed( -{ 2'b0,x177 }<<<3'd1 )+$signed( { 2'b0,x178 } <<<3'd1 )+$signed( { 2'b0,x179 } <<<3'd1 )+$signed( { 1'b0,x180 }  )+$signed( -{ 4'b0, x181 }<<<3'd3 )+$signed( -{ 1'b0,x182 } )+$signed( -{ 3'b0,x183 }<<<3'd2)+$signed( { 2'b0,x184 } <<<3'd1 )+$signed( -{ 3'b0,x185 }<<<3'd2)+$signed( { 2'b0,x186 } <<<3'd1 )+$signed( { 1'b0,x188 }  )+$signed( -{ 2'b0,x189 }<<<3'd1 )+$signed( { 1'b0,x190 }  )+$signed( { 3'b0,x191 }<<<3'd2 )+$signed( -{ 3'b0,x192 }<<<3'd2)+$signed( -{ 1'b0,x193 } )+$signed( -{ 2'b0,x194 }<<<3'd1 )+$signed( { 2'b0,x195 } <<<3'd1 )+$signed( { 2'b0,x196 } <<<3'd1 )+$signed( { 2'b0,x197 } <<<3'd1 )+$signed( -{ 2'b0,x198 }<<<3'd1 )+$signed( -{ 2'b0,x200 }<<<3'd1 )+$signed( -{ 2'b0,x202 }<<<3'd1 )+$signed( { 3'b0,x203 }<<<3'd2 )+$signed( { 2'b0,x204 } <<<3'd1 )+$signed( -{ 2'b0,x205 }<<<3'd1 )+$signed( { 1'b0,x206 }  )+$signed( { 3'b0,x208 }<<<3'd2 )+$signed( { 3'b0,x209 }<<<3'd2 )+$signed( { 1'b0,x210 }  )+$signed( { 1'b0,x211 }  )+$signed( -{ 1'b0,x213 } )+$signed( { 3'b0,x214 }<<<3'd2 )+$signed( { 1'b0,x215 }  )+$signed( { 2'b0,x216 } <<<3'd1 )+$signed( -{ 2'b0,x217 }<<<3'd1 )+$signed( { 2'b0,x218 } <<<3'd1 )+$signed( -{ 3'b0,x220 }<<<3'd2)+$signed( -{ 2'b0,x221 }<<<3'd1 )+$signed( -{ 2'b0,x222 }<<<3'd1 )+$signed( -{ 1'b0,x223 } )+$signed( { 2'b0,x224 } <<<3'd1 )+$signed( -{ 5'b0,x225 }<<<3'd4 )+$signed( { 2'b0,x226 } <<<3'd1 )+$signed( { 3'b0,x227 }<<<3'd2 )+$signed( -{ 2'b0,x228 }<<<3'd1 )+$signed( -{ 2'b0,x229 }<<<3'd1 )+$signed( -{ 1'b0,x230 } )+$signed( -{ 1'b0,x233 } )+$signed( { 3'b0,x235 }<<<3'd2 )+$signed( { 3'b0,x236 }<<<3'd2 )+$signed( -{ 1'b0,x237 } )+$signed( -{ 1'b0,x238 } )+$signed( -{ 1'b0,x239 } )+$signed( -{ 2'b0,x240 }<<<3'd1 )+$signed( -{ 1'b0,x241 } )+$signed( -{ 3'b0,x242 }<<<3'd2)+$signed( -{ 3'b0,x243 }<<<3'd2)+$signed( { 2'b0,x244 } <<<3'd1 )+$signed( { 3'b0,x245 }<<<3'd2 )+$signed( -{ 1'b0,x246 } )+$signed( -{ 2'b0,x247 }<<<3'd1 )+$signed( -{ 3'b0,x248 }<<<3'd2)+$signed( { 1'b0,x249 }  )+$signed( -{ 1'b0,x250 } )+$signed( -{ 1'b0,x251 } )+$signed( { 1'b0,x252 }  )+$signed( { 3'b0,x253 }<<<3'd2 )+$signed( { 2'b0,x254 } <<<3'd1 )+$signed( -{ 2'b0,x255 }<<<3'd1 )+$signed( -{ 2'b0,x256 }<<<3'd1 )+$signed( { 1'b0,x257 }  )+$signed( -{ 3'b0,x258 }<<<3'd2)+$signed( -{ 1'b0,x259 } )+$signed( -{ 1'b0,x260 } )+$signed( -{ 3'b0,x261 }<<<3'd2)+$signed( -{ 2'b0,x262 }<<<3'd1 )+$signed( { 3'b0,x263 }<<<3'd2 )+$signed( { 2'b0,x264 } <<<3'd1 )+$signed( { 1'b0,x265 }  )+$signed( { 3'b0,x267 }<<<3'd2 )+$signed( -{ 2'b0,x268 }<<<3'd1 )+$signed( { 2'b0,x269 } <<<3'd1 )+$signed( -{ 1'b0,x270 } )+$signed( { 1'b0,x271 }  )+$signed( -{ 3'b0,x272 }<<<3'd2)+$signed( -{ 1'b0,x273 } )+$signed( -{ 3'b0,x274 }<<<3'd2)+$signed( { 1'b0,x276 }  )+$signed( { 3'b0,x278 }<<<3'd2 )+$signed( -{ 4'b0, x279 }<<<3'd3 )+$signed( { 1'b0,x280 }  )+$signed( { 3'b0,x281 }<<<3'd2 )+$signed( -{ 1'b0,x284 } )+$signed( -{ 1'b0,x286 } )+$signed( -{ 3'b0,x288 }<<<3'd2)+$signed( { 3'b0,x289 }<<<3'd2 )+$signed( -{ 2'b0,x290 }<<<3'd1 )+$signed( { 1'b0,x291 }  )+$signed( -{ 3'b0,x292 }<<<3'd2)+$signed( -{ 2'b0,x293 }<<<3'd1 )+$signed( { 1'b0,x294 }  )+$signed( { 3'b0,x295 }<<<3'd2 )+$signed( -{ 3'b0,x296 }<<<3'd2)+$signed( -{ 3'b0,x299 }<<<3'd2)+$signed( { 1'b0,x300 }  )+$signed( -{ 3'b0,x301 }<<<3'd2)+$signed( -{ 2'b0,x302 }<<<3'd1 )+$signed( { 1'b0,x304 }  )+$signed( -{ 4'b0, x305 }<<<3'd3 )+$signed( -{ 3'b0,x306 }<<<3'd2)+$signed( -{ 3'b0,x307 }<<<3'd2)+$signed( -{ 1'b0,x308 } )+$signed( -{ 1'b0,x310 } )+$signed( -{ 3'b0,x312 }<<<3'd2)+$signed( { 1'b0,x313 }  )+$signed( { 1'b0,x314 }  )+$signed( { 2'b0,x315 } <<<3'd1 )+$signed( { 3'b0,x316 }<<<3'd2 )+$signed( -{ 1'b0,x317 } )+$signed( -{ 5'b0,x318 }<<<3'd4 )+$signed( -{ 2'b0,x319 }<<<3'd1 )+$signed( { 2'b0,x320 } <<<3'd1 )+$signed( { 3'b0,x321 }<<<3'd2 )+$signed( { 3'b0,x322 }<<<3'd2 )+$signed( -{ 3'b0,x323 }<<<3'd2)+$signed( -{ 1'b0,x326 } )+$signed( -{ 2'b0,x327 }<<<3'd1 )+$signed( { 3'b0,x328 }<<<3'd2 )+$signed( { 1'b0,x329 }  )+$signed( -{ 3'b0,x330 }<<<3'd2)+$signed( -{ 3'b0,x331 }<<<3'd2)+$signed( { 2'b0,x332 } <<<3'd1 )+$signed( { 3'b0,x333 }<<<3'd2 )+$signed( { 3'b0,x334 }<<<3'd2 )+$signed( -{ 1'b0,x335 } )+$signed( -{ 1'b0,x336 } )+$signed( -{ 3'b0,x338 }<<<3'd2)+$signed( -{ 2'b0,x339 }<<<3'd1 )+$signed( -{ 1'b0,x340 } )+$signed( { 3'b0,x341 }<<<3'd2 )+$signed( -{ 2'b0,x342 }<<<3'd1 )+$signed( { 3'b0,x343 }<<<3'd2 )+$signed( -{ 3'b0,x344 }<<<3'd2)+$signed( { 3'b0,x345 }<<<3'd2 )+$signed( { 2'b0,x346 } <<<3'd1 )+$signed( { 4'b0,x347 }<<<3'd3 )+$signed( -{ 2'b0,x348 }<<<3'd1 )+$signed( -{ 2'b0,x349 }<<<3'd1 )+$signed( -{ 1'b0,x350 } )+$signed( { 1'b0,x351 }  )+$signed( { 1'b0,x352 }  )+$signed( -{ 1'b0,x354 } )+$signed( { 2'b0,x355 } <<<3'd1 )+$signed( -{ 2'b0,x356 }<<<3'd1 )+$signed( { 3'b0,x357 }<<<3'd2 )+$signed( { 2'b0,x358 } <<<3'd1 )+$signed( -{ 3'b0,x359 }<<<3'd2)+$signed( { 2'b0,x360 } <<<3'd1 )+$signed( -{ 2'b0,x361 }<<<3'd1 )+$signed( { 2'b0,x362 } <<<3'd1 )+$signed( { 3'b0,x363 }<<<3'd2 )+$signed( { 3'b0,x364 }<<<3'd2 )+$signed( -{ 2'b0,x365 }<<<3'd1 )+$signed( -{ 3'b0,x366 }<<<3'd2)+$signed( -{ 2'b0,x367 }<<<3'd1 )+$signed( { 1'b0,x368 }  )+$signed( -{ 4'b0, x369 }<<<3'd3 )+$signed( -{ 2'b0,x370 }<<<3'd1 )+$signed( { 2'b0,x371 } <<<3'd1 )+$signed( -{ 1'b0,x372 } )+$signed( { 2'b0,x373 } <<<3'd1 )+$signed( -{ 2'b0,x374 }<<<3'd1 )+$signed( { 1'b0,x375 }  )+$signed( -{ 1'b0,x376 } )+$signed( -{ 3'b0,x377 }<<<3'd2)+$signed( -{ 3'b0,x378 }<<<3'd2)+$signed( { 1'b0,x380 }  )+$signed( -{ 3'b0,x381 }<<<3'd2)+$signed( -{ 2'b0,x382 }<<<3'd1 )+$signed( -{ 3'b0,x383 }<<<3'd2)+$signed( { 3'b0,x384 }<<<3'd2 )+$signed( { 1'b0,x385 }  )+$signed( { 3'b0,x386 }<<<3'd2 )+$signed( { 3'b0,x387 }<<<3'd2 )+$signed( -{ 3'b0,x388 }<<<3'd2)+$signed( { 1'b0,x389 }  )+$signed( -{ 3'b0,x390 }<<<3'd2)+$signed( -{ 2'b0,x391 }<<<3'd1 )+$signed( -{ 2'b0,x392 }<<<3'd1 )+$signed( { 3'b0,x393 }<<<3'd2 )+$signed( -{ 3'b0,x394 }<<<3'd2)+$signed( -{ 1'b0,x395 } )+$signed( -{ 3'b0,x396 }<<<3'd2)+$signed( -{ 2'b0,x397 }<<<3'd1 )+$signed( -{ 2'b0,x398 }<<<3'd1 )+$signed( { 3'b0,x399 }<<<3'd2 )+$signed( { 2'b0,x401 } <<<3'd1 )+$signed( -{ 3'b0,x402 }<<<3'd2)+$signed( -{ 4'b0, x403 }<<<3'd3 )+$signed( -{ 2'b0,x404 }<<<3'd1 )+$signed( -{ 3'b0,x405 }<<<3'd2)+$signed( { 2'b0,x406 } <<<3'd1 )+$signed( -{ 3'b0,x407 }<<<3'd2)+$signed( { 2'b0,x408 } <<<3'd1 )+$signed( { 3'b0,x409 }<<<3'd2 )+$signed( { 2'b0,x410 } <<<3'd1 )+$signed( { 2'b0,x412 } <<<3'd1 )+$signed( { 1'b0,x413 }  )+$signed( { 1'b0,x414 }  )+$signed( { 2'b0,x415 } <<<3'd1 )+$signed( -{ 3'b0,x416 }<<<3'd2)+$signed( -{ 3'b0,x417 }<<<3'd2)+$signed( -{ 1'b0,x418 } )+$signed( { 1'b0,x419 }  )+$signed( -{ 3'b0,x420 }<<<3'd2)+$signed( -{ 1'b0,x422 } )+$signed( { 2'b0,x423 } <<<3'd1 )+$signed( { 1'b0,x424 }  )+$signed( { 3'b0,x425 }<<<3'd2 )+$signed( -{ 1'b0,x426 } )+$signed( { 1'b0,x427 }  )+$signed( -{ 1'b0,x429 } )+$signed( -{ 3'b0,x430 }<<<3'd2)+$signed( { 2'b0,x431 } <<<3'd1 )+$signed( -{ 1'b0,x432 } )+$signed( { 2'b0,x433 } <<<3'd1 )+$signed( { 2'b0,x434 } <<<3'd1 )+$signed( -{ 4'b0, x435 }<<<3'd3 )+$signed( { 2'b0,x436 } <<<3'd1 )+$signed( -{ 2'b0,x437 }<<<3'd1 )+$signed( { 2'b0,x438 } <<<3'd1 )+$signed( -{ 3'b0,x439 }<<<3'd2)+$signed( -{ 3'b0,x440 }<<<3'd2)+$signed( -{ 1'b0,x441 } )+$signed( { 3'b0,x442 }<<<3'd2 )+$signed( -{ 3'b0,x443 }<<<3'd2)+$signed( -{ 2'b0,x444 }<<<3'd1 )+$signed( -{ 1'b0,x445 } )+$signed( -{ 3'b0,x446 }<<<3'd2)+$signed( { 2'b0,x447 } <<<3'd1 )+$signed( -{ 3'b0,x448 }<<<3'd2)+$signed( -{ 2'b0,x450 }<<<3'd1 )+$signed( -{ 1'b0,x451 } )+$signed( { 2'b0,x452 } <<<3'd1 )+$signed( { 2'b0,x453 } <<<3'd1 )+$signed( -{ 1'b0,x455 } )+$signed( -{ 3'b0,x456 }<<<3'd2)+$signed( -{ 2'b0,x457 }<<<3'd1 )+$signed( { 1'b0,x458 }  )+$signed( -{ 2'b0,x459 }<<<3'd1 )+$signed( { 3'b0,x460 }<<<3'd2 )+$signed( -{ 3'b0,x461 }<<<3'd2)+$signed( { 2'b0,x462 } <<<3'd1 )+$signed( { 3'b0,x463 }<<<3'd2 )+$signed( { 2'b0,x464 } <<<3'd1 )+$signed( { 3'b0,x465 }<<<3'd2 )+$signed( { 2'b0,x466 } <<<3'd1 )+$signed( { 3'b0,x468 }<<<3'd2 )+$signed( -{ 4'b0, x469 }<<<3'd3 )+$signed( { 1'b0,x470 }  )+$signed( { 4'b0,x471 }<<<3'd3 )+$signed( -{ 2'b0,x472 }<<<3'd1 )+$signed( { 3'b0,x473 }<<<3'd2 )+$signed( -{ 3'b0,x474 }<<<3'd2)+$signed( { 2'b0,x476 } <<<3'd1 )+$signed( { 2'b0,x477 } <<<3'd1 )+$signed( -{ 1'b0,x479 } )+$signed( { 3'b0,x480 }<<<3'd2 )+$signed( -{ 3'b0,x481 }<<<3'd2)+$signed( -{ 3'b0,x482 }<<<3'd2)+$signed( { 2'b0,x483 } <<<3'd1 )+$signed( { 3'b0,x484 }<<<3'd2 )+$signed( -{ 2'b0,x485 }<<<3'd1 )+$signed( { 2'b0,x486 } <<<3'd1 )+$signed( -{ 2'b0,x487 }<<<3'd1 )+$signed( { 1'b0,x488 }  )+$signed( -{ 2'b0,x489 }<<<3'd1 )+$signed( { 3'b0,x490 }<<<3'd2 )+$signed( -{ 3'b0,x491 }<<<3'd2)+$signed( -{ 1'b0,x492 } )+$signed( { 2'b0,x493 } <<<3'd1 )+$signed( -{ 3'b0,x494 }<<<3'd2)+$signed( -{ 4'b0, x495 }<<<3'd3 )+$signed(13'd56);
assign y15=temp_y[15][13] ==1'b1 ? 6'd0 :  
    temp_y[15][10] ==1'b1 ? 6'd63 : 
    temp_y[15][3]==1'b1 ? temp_y[15][9:4]+1'b1 : temp_y[15][9:4];
assign temp_y[16] = 
+$signed( { 1'b0,x0 }  )+$signed( { 1'b0,x1 }  )+$signed( -{ 1'b0,x2 } )+$signed( -{ 3'b0,x3 }<<<3'd2)+$signed( -{ 1'b0,x4 } )+$signed( -{ 1'b0,x5 } )+$signed( { 1'b0,x6 }  )+$signed( { 2'b0,x7 } <<<3'd1 )+$signed( { 2'b0,x8 } <<<3'd1 )+$signed( -{ 3'b0,x9 }<<<3'd2)+$signed( { 2'b0,x10 } <<<3'd1 )+$signed( { 1'b0,x11 }  )+$signed( -{ 2'b0,x12 }<<<3'd1 )+$signed( { 3'b0,x13 }<<<3'd2 )+$signed( { 3'b0,x15 }<<<3'd2 )+$signed( -{ 1'b0,x16 } )+$signed( -{ 4'b0, x17 }<<<3'd3 )+$signed( -{ 1'b0,x19 } )+$signed( -{ 1'b0,x20 } )+$signed( -{ 2'b0,x21 }<<<3'd1 )+$signed( -{ 1'b0,x22 } )+$signed( -{ 2'b0,x23 }<<<3'd1 )+$signed( { 2'b0,x24 } <<<3'd1 )+$signed( { 3'b0,x25 }<<<3'd2 )+$signed( -{ 3'b0,x26 }<<<3'd2)+$signed( { 1'b0,x28 }  )+$signed( -{ 3'b0,x29 }<<<3'd2)+$signed( -{ 3'b0,x30 }<<<3'd2)+$signed( -{ 1'b0,x31 } )+$signed( { 2'b0,x32 } <<<3'd1 )+$signed( { 2'b0,x33 } <<<3'd1 )+$signed( { 1'b0,x34 }  )+$signed( -{ 2'b0,x35 }<<<3'd1 )+$signed( { 2'b0,x36 } <<<3'd1 )+$signed( { 3'b0,x37 }<<<3'd2 )+$signed( { 1'b0,x38 }  )+$signed( { 1'b0,x40 }  )+$signed( -{ 3'b0,x41 }<<<3'd2)+$signed( { 3'b0,x42 }<<<3'd2 )+$signed( -{ 1'b0,x43 } )+$signed( -{ 2'b0,x44 }<<<3'd1 )+$signed( { 3'b0,x45 }<<<3'd2 )+$signed( -{ 1'b0,x47 } )+$signed( { 2'b0,x48 } <<<3'd1 )+$signed( { 1'b0,x49 }  )+$signed( -{ 2'b0,x50 }<<<3'd1 )+$signed( { 2'b0,x52 } <<<3'd1 )+$signed( -{ 4'b0, x53 }<<<3'd3 )+$signed( -{ 2'b0,x54 }<<<3'd1 )+$signed( { 3'b0,x55 }<<<3'd2 )+$signed( { 2'b0,x56 } <<<3'd1 )+$signed( { 2'b0,x57 } <<<3'd1 )+$signed( -{ 3'b0,x58 }<<<3'd2)+$signed( -{ 3'b0,x59 }<<<3'd2)+$signed( { 2'b0,x60 } <<<3'd1 )+$signed( { 3'b0,x61 }<<<3'd2 )+$signed( { 2'b0,x62 } <<<3'd1 )+$signed( -{ 4'b0, x63 }<<<3'd3 )+$signed( -{ 3'b0,x64 }<<<3'd2)+$signed( -{ 3'b0,x65 }<<<3'd2)+$signed( { 3'b0,x66 }<<<3'd2 )+$signed( -{ 1'b0,x67 } )+$signed( -{ 3'b0,x68 }<<<3'd2)+$signed( -{ 2'b0,x70 }<<<3'd1 )+$signed( -{ 3'b0,x71 }<<<3'd2)+$signed( { 1'b0,x72 }  )+$signed( { 2'b0,x73 } <<<3'd1 )+$signed( { 2'b0,x74 } <<<3'd1 )+$signed( -{ 3'b0,x75 }<<<3'd2)+$signed( { 3'b0,x76 }<<<3'd2 )+$signed( -{ 3'b0,x77 }<<<3'd2)+$signed( { 3'b0,x79 }<<<3'd2 )+$signed( { 1'b0,x80 }  )+$signed( -{ 2'b0,x81 }<<<3'd1 )+$signed( { 1'b0,x82 }  )+$signed( { 2'b0,x83 } <<<3'd1 )+$signed( { 1'b0,x84 }  )+$signed( { 2'b0,x85 } <<<3'd1 )+$signed( { 3'b0,x86 }<<<3'd2 )+$signed( { 2'b0,x87 } <<<3'd1 )+$signed( -{ 2'b0,x88 }<<<3'd1 )+$signed( -{ 4'b0, x89 }<<<3'd3 )+$signed( -{ 2'b0,x90 }<<<3'd1 )+$signed( { 2'b0,x91 } <<<3'd1 )+$signed( -{ 2'b0,x93 }<<<3'd1 )+$signed( -{ 1'b0,x95 } )+$signed( -{ 3'b0,x96 }<<<3'd2)+$signed( { 1'b0,x97 }  )+$signed( -{ 3'b0,x98 }<<<3'd2)+$signed( { 3'b0,x99 }<<<3'd2 )+$signed( { 3'b0,x100 }<<<3'd2 )+$signed( { 1'b0,x101 }  )+$signed( { 4'b0,x102 }<<<3'd3 )+$signed( { 4'b0,x104 }<<<3'd3 )+$signed( { 3'b0,x105 }<<<3'd2 )+$signed( { 2'b0,x106 } <<<3'd1 )+$signed( { 3'b0,x107 }<<<3'd2 )+$signed( -{ 1'b0,x108 } )+$signed( { 1'b0,x110 }  )+$signed( -{ 4'b0, x111 }<<<3'd3 )+$signed( { 3'b0,x112 }<<<3'd2 )+$signed( { 3'b0,x113 }<<<3'd2 )+$signed( -{ 3'b0,x114 }<<<3'd2)+$signed( { 3'b0,x115 }<<<3'd2 )+$signed( -{ 3'b0,x116 }<<<3'd2)+$signed( { 4'b0,x117 }<<<3'd3 )+$signed( { 4'b0,x118 }<<<3'd3 )+$signed( { 1'b0,x119 }  )+$signed( { 4'b0,x120 }<<<3'd3 )+$signed( { 3'b0,x121 }<<<3'd2 )+$signed( { 3'b0,x122 }<<<3'd2 )+$signed( -{ 1'b0,x123 } )+$signed( { 1'b0,x124 }  )+$signed( -{ 2'b0,x125 }<<<3'd1 )+$signed( -{ 1'b0,x126 } )+$signed( -{ 2'b0,x127 }<<<3'd1 )+$signed( -{ 1'b0,x128 } )+$signed( -{ 4'b0, x129 }<<<3'd3 )+$signed( -{ 2'b0,x130 }<<<3'd1 )+$signed( -{ 3'b0,x131 }<<<3'd2)+$signed( { 2'b0,x132 } <<<3'd1 )+$signed( -{ 3'b0,x133 }<<<3'd2)+$signed( -{ 4'b0, x135 }<<<3'd3 )+$signed( -{ 2'b0,x136 }<<<3'd1 )+$signed( -{ 3'b0,x137 }<<<3'd2)+$signed( { 4'b0,x138 }<<<3'd3 )+$signed( { 2'b0,x139 } <<<3'd1 )+$signed( { 3'b0,x140 }<<<3'd2 )+$signed( -{ 2'b0,x141 }<<<3'd1 )+$signed( { 2'b0,x142 } <<<3'd1 )+$signed( -{ 4'b0, x143 }<<<3'd3 )+$signed( -{ 3'b0,x144 }<<<3'd2)+$signed( -{ 1'b0,x145 } )+$signed( { 2'b0,x146 } <<<3'd1 )+$signed( { 1'b0,x147 }  )+$signed( { 2'b0,x148 } <<<3'd1 )+$signed( { 3'b0,x150 }<<<3'd2 )+$signed( -{ 2'b0,x151 }<<<3'd1 )+$signed( { 2'b0,x152 } <<<3'd1 )+$signed( -{ 3'b0,x153 }<<<3'd2)+$signed( -{ 3'b0,x154 }<<<3'd2)+$signed( -{ 3'b0,x156 }<<<3'd2)+$signed( { 1'b0,x157 }  )+$signed( { 4'b0,x158 }<<<3'd3 )+$signed( { 3'b0,x159 }<<<3'd2 )+$signed( -{ 4'b0, x161 }<<<3'd3 )+$signed( { 3'b0,x163 }<<<3'd2 )+$signed( { 3'b0,x165 }<<<3'd2 )+$signed( { 3'b0,x166 }<<<3'd2 )+$signed( { 2'b0,x167 } <<<3'd1 )+$signed( -{ 3'b0,x168 }<<<3'd2)+$signed( { 3'b0,x169 }<<<3'd2 )+$signed( { 3'b0,x171 }<<<3'd2 )+$signed( { 3'b0,x172 }<<<3'd2 )+$signed( -{ 1'b0,x173 } )+$signed( { 3'b0,x174 }<<<3'd2 )+$signed( -{ 2'b0,x175 }<<<3'd1 )+$signed( -{ 1'b0,x176 } )+$signed( { 1'b0,x177 }  )+$signed( -{ 2'b0,x178 }<<<3'd1 )+$signed( -{ 2'b0,x179 }<<<3'd1 )+$signed( { 2'b0,x180 } <<<3'd1 )+$signed( { 3'b0,x181 }<<<3'd2 )+$signed( -{ 2'b0,x182 }<<<3'd1 )+$signed( { 3'b0,x183 }<<<3'd2 )+$signed( { 3'b0,x184 }<<<3'd2 )+$signed( -{ 2'b0,x185 }<<<3'd1 )+$signed( -{ 3'b0,x186 }<<<3'd2)+$signed( { 1'b0,x187 }  )+$signed( { 1'b0,x188 }  )+$signed( -{ 1'b0,x189 } )+$signed( { 2'b0,x190 } <<<3'd1 )+$signed( { 1'b0,x191 }  )+$signed( { 1'b0,x192 }  )+$signed( -{ 3'b0,x193 }<<<3'd2)+$signed( { 1'b0,x194 }  )+$signed( -{ 3'b0,x196 }<<<3'd2)+$signed( { 1'b0,x197 }  )+$signed( -{ 2'b0,x198 }<<<3'd1 )+$signed( -{ 2'b0,x199 }<<<3'd1 )+$signed( -{ 2'b0,x200 }<<<3'd1 )+$signed( { 3'b0,x201 }<<<3'd2 )+$signed( -{ 3'b0,x202 }<<<3'd2)+$signed( -{ 3'b0,x203 }<<<3'd2)+$signed( { 3'b0,x205 }<<<3'd2 )+$signed( { 2'b0,x206 } <<<3'd1 )+$signed( { 2'b0,x207 } <<<3'd1 )+$signed( { 2'b0,x208 } <<<3'd1 )+$signed( -{ 2'b0,x209 }<<<3'd1 )+$signed( { 2'b0,x210 } <<<3'd1 )+$signed( -{ 2'b0,x211 }<<<3'd1 )+$signed( -{ 2'b0,x212 }<<<3'd1 )+$signed( -{ 2'b0,x213 }<<<3'd1 )+$signed( { 3'b0,x214 }<<<3'd2 )+$signed( -{ 3'b0,x215 }<<<3'd2)+$signed( -{ 1'b0,x216 } )+$signed( -{ 3'b0,x217 }<<<3'd2)+$signed( { 1'b0,x218 }  )+$signed( { 1'b0,x219 }  )+$signed( -{ 4'b0, x221 }<<<3'd3 )+$signed( -{ 3'b0,x222 }<<<3'd2)+$signed( { 2'b0,x223 } <<<3'd1 )+$signed( -{ 2'b0,x224 }<<<3'd1 )+$signed( { 3'b0,x225 }<<<3'd2 )+$signed( -{ 3'b0,x226 }<<<3'd2)+$signed( -{ 2'b0,x227 }<<<3'd1 )+$signed( -{ 2'b0,x228 }<<<3'd1 )+$signed( -{ 3'b0,x229 }<<<3'd2)+$signed( -{ 4'b0, x230 }<<<3'd3 )+$signed( { 2'b0,x231 } <<<3'd1 )+$signed( -{ 1'b0,x232 } )+$signed( -{ 3'b0,x233 }<<<3'd2)+$signed( { 3'b0,x234 }<<<3'd2 )+$signed( { 1'b0,x235 }  )+$signed( { 3'b0,x236 }<<<3'd2 )+$signed( -{ 2'b0,x237 }<<<3'd1 )+$signed( { 3'b0,x238 }<<<3'd2 )+$signed( -{ 1'b0,x239 } )+$signed( -{ 3'b0,x241 }<<<3'd2)+$signed( -{ 2'b0,x242 }<<<3'd1 )+$signed( { 2'b0,x243 } <<<3'd1 )+$signed( -{ 3'b0,x244 }<<<3'd2)+$signed( { 2'b0,x245 } <<<3'd1 )+$signed( -{ 1'b0,x246 } )+$signed( -{ 3'b0,x247 }<<<3'd2)+$signed( -{ 1'b0,x248 } )+$signed( { 3'b0,x249 }<<<3'd2 )+$signed( -{ 3'b0,x250 }<<<3'd2)+$signed( -{ 3'b0,x251 }<<<3'd2)+$signed( { 1'b0,x252 }  )+$signed( { 4'b0,x253 }<<<3'd3 )+$signed( -{ 4'b0, x254 }<<<3'd3 )+$signed( -{ 1'b0,x255 } )+$signed( { 2'b0,x256 } <<<3'd1 )+$signed( -{ 3'b0,x258 }<<<3'd2)+$signed( -{ 2'b0,x260 }<<<3'd1 )+$signed( -{ 1'b0,x261 } )+$signed( -{ 3'b0,x262 }<<<3'd2)+$signed( { 1'b0,x263 }  )+$signed( -{ 2'b0,x264 }<<<3'd1 )+$signed( -{ 2'b0,x266 }<<<3'd1 )+$signed( { 1'b0,x267 }  )+$signed( { 1'b0,x269 }  )+$signed( { 2'b0,x270 } <<<3'd1 )+$signed( -{ 5'b0,x271 }<<<3'd4 )+$signed( -{ 1'b0,x272 } )+$signed( { 1'b0,x273 }  )+$signed( -{ 1'b0,x274 } )+$signed( -{ 2'b0,x275 }<<<3'd1 )+$signed( -{ 1'b0,x276 } )+$signed( { 3'b0,x277 }<<<3'd2 )+$signed( -{ 2'b0,x279 }<<<3'd1 )+$signed( { 1'b0,x280 }  )+$signed( -{ 3'b0,x281 }<<<3'd2)+$signed( -{ 2'b0,x282 }<<<3'd1 )+$signed( -{ 2'b0,x284 }<<<3'd1 )+$signed( -{ 1'b0,x285 } )+$signed( -{ 1'b0,x286 } )+$signed( -{ 3'b0,x287 }<<<3'd2)+$signed( -{ 2'b0,x288 }<<<3'd1 )+$signed( { 3'b0,x291 }<<<3'd2 )+$signed( { 2'b0,x292 } <<<3'd1 )+$signed( -{ 1'b0,x293 } )+$signed( { 2'b0,x295 } <<<3'd1 )+$signed( -{ 1'b0,x296 } )+$signed( { 2'b0,x297 } <<<3'd1 )+$signed( { 3'b0,x298 }<<<3'd2 )+$signed( -{ 3'b0,x299 }<<<3'd2)+$signed( { 3'b0,x300 }<<<3'd2 )+$signed( { 3'b0,x301 }<<<3'd2 )+$signed( -{ 3'b0,x302 }<<<3'd2)+$signed( { 2'b0,x303 } <<<3'd1 )+$signed( { 2'b0,x304 } <<<3'd1 )+$signed( -{ 2'b0,x305 }<<<3'd1 )+$signed( -{ 1'b0,x306 } )+$signed( { 1'b0,x307 }  )+$signed( { 2'b0,x308 } <<<3'd1 )+$signed( { 1'b0,x309 }  )+$signed( -{ 3'b0,x310 }<<<3'd2)+$signed( { 4'b0,x311 }<<<3'd3 )+$signed( -{ 2'b0,x312 }<<<3'd1 )+$signed( { 2'b0,x313 } <<<3'd1 )+$signed( { 1'b0,x314 }  )+$signed( -{ 3'b0,x315 }<<<3'd2)+$signed( -{ 3'b0,x316 }<<<3'd2)+$signed( { 3'b0,x317 }<<<3'd2 )+$signed( { 3'b0,x318 }<<<3'd2 )+$signed( -{ 3'b0,x319 }<<<3'd2)+$signed( { 2'b0,x320 } <<<3'd1 )+$signed( -{ 2'b0,x321 }<<<3'd1 )+$signed( -{ 3'b0,x322 }<<<3'd2)+$signed( { 1'b0,x323 }  )+$signed( { 1'b0,x324 }  )+$signed( -{ 4'b0, x325 }<<<3'd3 )+$signed( { 1'b0,x326 }  )+$signed( -{ 2'b0,x328 }<<<3'd1 )+$signed( -{ 1'b0,x329 } )+$signed( { 3'b0,x330 }<<<3'd2 )+$signed( { 3'b0,x331 }<<<3'd2 )+$signed( -{ 1'b0,x332 } )+$signed( { 3'b0,x333 }<<<3'd2 )+$signed( -{ 2'b0,x334 }<<<3'd1 )+$signed( -{ 1'b0,x335 } )+$signed( { 1'b0,x336 }  )+$signed( -{ 4'b0, x338 }<<<3'd3 )+$signed( { 3'b0,x339 }<<<3'd2 )+$signed( { 3'b0,x340 }<<<3'd2 )+$signed( -{ 3'b0,x341 }<<<3'd2)+$signed( -{ 1'b0,x342 } )+$signed( { 2'b0,x343 } <<<3'd1 )+$signed( { 3'b0,x344 }<<<3'd2 )+$signed( { 1'b0,x345 }  )+$signed( -{ 3'b0,x347 }<<<3'd2)+$signed( -{ 2'b0,x348 }<<<3'd1 )+$signed( { 1'b0,x349 }  )+$signed( { 1'b0,x350 }  )+$signed( -{ 3'b0,x351 }<<<3'd2)+$signed( -{ 2'b0,x352 }<<<3'd1 )+$signed( -{ 3'b0,x353 }<<<3'd2)+$signed( { 1'b0,x354 }  )+$signed( -{ 4'b0, x355 }<<<3'd3 )+$signed( { 2'b0,x356 } <<<3'd1 )+$signed( { 3'b0,x357 }<<<3'd2 )+$signed( { 2'b0,x358 } <<<3'd1 )+$signed( -{ 1'b0,x359 } )+$signed( -{ 3'b0,x360 }<<<3'd2)+$signed( { 2'b0,x361 } <<<3'd1 )+$signed( { 4'b0,x362 }<<<3'd3 )+$signed( -{ 3'b0,x363 }<<<3'd2)+$signed( -{ 5'b0,x364 }<<<3'd4 )+$signed( { 3'b0,x365 }<<<3'd2 )+$signed( -{ 3'b0,x366 }<<<3'd2)+$signed( { 3'b0,x367 }<<<3'd2 )+$signed( -{ 2'b0,x368 }<<<3'd1 )+$signed( -{ 1'b0,x370 } )+$signed( { 3'b0,x371 }<<<3'd2 )+$signed( { 1'b0,x372 }  )+$signed( { 2'b0,x373 } <<<3'd1 )+$signed( -{ 2'b0,x374 }<<<3'd1 )+$signed( -{ 2'b0,x375 }<<<3'd1 )+$signed( -{ 2'b0,x376 }<<<3'd1 )+$signed( -{ 2'b0,x377 }<<<3'd1 )+$signed( { 3'b0,x378 }<<<3'd2 )+$signed( -{ 2'b0,x379 }<<<3'd1 )+$signed( -{ 1'b0,x380 } )+$signed( -{ 3'b0,x381 }<<<3'd2)+$signed( { 2'b0,x382 } <<<3'd1 )+$signed( -{ 3'b0,x383 }<<<3'd2)+$signed( { 3'b0,x384 }<<<3'd2 )+$signed( { 3'b0,x385 }<<<3'd2 )+$signed( -{ 3'b0,x387 }<<<3'd2)+$signed( { 2'b0,x388 } <<<3'd1 )+$signed( -{ 2'b0,x389 }<<<3'd1 )+$signed( { 3'b0,x390 }<<<3'd2 )+$signed( -{ 2'b0,x391 }<<<3'd1 )+$signed( { 3'b0,x392 }<<<3'd2 )+$signed( -{ 3'b0,x393 }<<<3'd2)+$signed( -{ 3'b0,x394 }<<<3'd2)+$signed( -{ 3'b0,x395 }<<<3'd2)+$signed( -{ 2'b0,x396 }<<<3'd1 )+$signed( -{ 3'b0,x397 }<<<3'd2)+$signed( { 3'b0,x398 }<<<3'd2 )+$signed( { 1'b0,x399 }  )+$signed( { 4'b0,x400 }<<<3'd3 )+$signed( { 3'b0,x401 }<<<3'd2 )+$signed( { 3'b0,x403 }<<<3'd2 )+$signed( -{ 2'b0,x404 }<<<3'd1 )+$signed( { 2'b0,x405 } <<<3'd1 )+$signed( -{ 2'b0,x406 }<<<3'd1 )+$signed( { 1'b0,x407 }  )+$signed( { 3'b0,x408 }<<<3'd2 )+$signed( -{ 1'b0,x409 } )+$signed( -{ 3'b0,x410 }<<<3'd2)+$signed( { 3'b0,x411 }<<<3'd2 )+$signed( -{ 3'b0,x412 }<<<3'd2)+$signed( { 3'b0,x413 }<<<3'd2 )+$signed( -{ 3'b0,x414 }<<<3'd2)+$signed( -{ 2'b0,x415 }<<<3'd1 )+$signed( { 3'b0,x416 }<<<3'd2 )+$signed( { 3'b0,x417 }<<<3'd2 )+$signed( { 3'b0,x418 }<<<3'd2 )+$signed( -{ 3'b0,x419 }<<<3'd2)+$signed( { 4'b0,x420 }<<<3'd3 )+$signed( -{ 3'b0,x421 }<<<3'd2)+$signed( -{ 3'b0,x422 }<<<3'd2)+$signed( -{ 2'b0,x423 }<<<3'd1 )+$signed( -{ 2'b0,x424 }<<<3'd1 )+$signed( -{ 2'b0,x425 }<<<3'd1 )+$signed( -{ 2'b0,x426 }<<<3'd1 )+$signed( { 2'b0,x427 } <<<3'd1 )+$signed( -{ 2'b0,x428 }<<<3'd1 )+$signed( { 3'b0,x429 }<<<3'd2 )+$signed( { 3'b0,x430 }<<<3'd2 )+$signed( { 3'b0,x431 }<<<3'd2 )+$signed( -{ 2'b0,x432 }<<<3'd1 )+$signed( { 2'b0,x433 } <<<3'd1 )+$signed( -{ 3'b0,x434 }<<<3'd2)+$signed( -{ 3'b0,x435 }<<<3'd2)+$signed( { 3'b0,x436 }<<<3'd2 )+$signed( { 2'b0,x437 } <<<3'd1 )+$signed( { 3'b0,x438 }<<<3'd2 )+$signed( { 3'b0,x439 }<<<3'd2 )+$signed( -{ 2'b0,x440 }<<<3'd1 )+$signed( { 2'b0,x441 } <<<3'd1 )+$signed( { 3'b0,x442 }<<<3'd2 )+$signed( -{ 3'b0,x444 }<<<3'd2)+$signed( -{ 2'b0,x445 }<<<3'd1 )+$signed( -{ 1'b0,x447 } )+$signed( -{ 3'b0,x448 }<<<3'd2)+$signed( -{ 4'b0, x449 }<<<3'd3 )+$signed( { 3'b0,x450 }<<<3'd2 )+$signed( -{ 2'b0,x451 }<<<3'd1 )+$signed( { 4'b0,x452 }<<<3'd3 )+$signed( -{ 2'b0,x453 }<<<3'd1 )+$signed( { 3'b0,x454 }<<<3'd2 )+$signed( { 3'b0,x455 }<<<3'd2 )+$signed( -{ 2'b0,x457 }<<<3'd1 )+$signed( -{ 2'b0,x458 }<<<3'd1 )+$signed( -{ 3'b0,x460 }<<<3'd2)+$signed( { 4'b0,x461 }<<<3'd3 )+$signed( -{ 3'b0,x462 }<<<3'd2)+$signed( { 2'b0,x463 } <<<3'd1 )+$signed( -{ 2'b0,x464 }<<<3'd1 )+$signed( -{ 4'b0, x466 }<<<3'd3 )+$signed( -{ 3'b0,x467 }<<<3'd2)+$signed( { 3'b0,x468 }<<<3'd2 )+$signed( { 3'b0,x469 }<<<3'd2 )+$signed( { 2'b0,x470 } <<<3'd1 )+$signed( -{ 1'b0,x471 } )+$signed( { 3'b0,x472 }<<<3'd2 )+$signed( { 2'b0,x473 } <<<3'd1 )+$signed( { 3'b0,x474 }<<<3'd2 )+$signed( { 2'b0,x475 } <<<3'd1 )+$signed( { 3'b0,x476 }<<<3'd2 )+$signed( -{ 3'b0,x477 }<<<3'd2)+$signed( { 1'b0,x478 }  )+$signed( { 2'b0,x479 } <<<3'd1 )+$signed( { 1'b0,x480 }  )+$signed( { 1'b0,x481 }  )+$signed( { 4'b0,x482 }<<<3'd3 )+$signed( { 3'b0,x483 }<<<3'd2 )+$signed( -{ 3'b0,x484 }<<<3'd2)+$signed( -{ 2'b0,x485 }<<<3'd1 )+$signed( -{ 3'b0,x488 }<<<3'd2)+$signed( { 2'b0,x489 } <<<3'd1 )+$signed( -{ 1'b0,x490 } )+$signed( -{ 3'b0,x491 }<<<3'd2)+$signed( { 3'b0,x493 }<<<3'd2 )+$signed( { 4'b0,x494 }<<<3'd3 )+$signed( { 2'b0,x495 } <<<3'd1 )-$signed(13'd0);
assign y16=temp_y[16][13] ==1'b1 ? 6'd0 :  
    temp_y[16][10] ==1'b1 ? 6'd63 : 
    temp_y[16][3]==1'b1 ? temp_y[16][9:4]+1'b1 : temp_y[16][9:4];
assign temp_y[17] = 
+$signed( -{ 3'b0,x0 }<<<3'd2)+$signed( { 1'b0,x1 }  )+$signed( { 2'b0,x2 } <<<3'd1 )+$signed( { 2'b0,x3 } <<<3'd1 )+$signed( { 3'b0,x4 }<<<3'd2 )+$signed( -{ 3'b0,x5 }<<<3'd2)+$signed( -{ 5'b0,x6 }<<<3'd4 )+$signed( { 1'b0,x7 }  )+$signed( -{ 3'b0,x8 }<<<3'd2)+$signed( { 1'b0,x9 }  )+$signed( { 2'b0,x10 } <<<3'd1 )+$signed( -{ 2'b0,x11 }<<<3'd1 )+$signed( { 3'b0,x12 }<<<3'd2 )+$signed( -{ 2'b0,x13 }<<<3'd1 )+$signed( { 3'b0,x14 }<<<3'd2 )+$signed( { 2'b0,x15 } <<<3'd1 )+$signed( { 1'b0,x16 }  )+$signed( -{ 3'b0,x17 }<<<3'd2)+$signed( -{ 2'b0,x18 }<<<3'd1 )+$signed( -{ 2'b0,x19 }<<<3'd1 )+$signed( { 1'b0,x20 }  )+$signed( { 2'b0,x21 } <<<3'd1 )+$signed( { 2'b0,x22 } <<<3'd1 )+$signed( -{ 3'b0,x23 }<<<3'd2)+$signed( { 3'b0,x24 }<<<3'd2 )+$signed( { 3'b0,x25 }<<<3'd2 )+$signed( -{ 2'b0,x26 }<<<3'd1 )+$signed( -{ 2'b0,x27 }<<<3'd1 )+$signed( { 1'b0,x28 }  )+$signed( -{ 2'b0,x29 }<<<3'd1 )+$signed( -{ 1'b0,x31 } )+$signed( { 3'b0,x32 }<<<3'd2 )+$signed( { 3'b0,x33 }<<<3'd2 )+$signed( { 2'b0,x34 } <<<3'd1 )+$signed( -{ 3'b0,x35 }<<<3'd2)+$signed( { 1'b0,x36 }  )+$signed( -{ 3'b0,x37 }<<<3'd2)+$signed( { 3'b0,x38 }<<<3'd2 )+$signed( { 3'b0,x39 }<<<3'd2 )+$signed( { 3'b0,x40 }<<<3'd2 )+$signed( -{ 3'b0,x41 }<<<3'd2)+$signed( -{ 4'b0, x42 }<<<3'd3 )+$signed( { 4'b0,x43 }<<<3'd3 )+$signed( { 3'b0,x44 }<<<3'd2 )+$signed( -{ 3'b0,x46 }<<<3'd2)+$signed( -{ 2'b0,x47 }<<<3'd1 )+$signed( -{ 5'b0,x48 }<<<3'd4 )+$signed( -{ 3'b0,x49 }<<<3'd2)+$signed( { 3'b0,x50 }<<<3'd2 )+$signed( -{ 2'b0,x51 }<<<3'd1 )+$signed( -{ 4'b0, x52 }<<<3'd3 )+$signed( -{ 1'b0,x53 } )+$signed( { 4'b0,x54 }<<<3'd3 )+$signed( -{ 3'b0,x55 }<<<3'd2)+$signed( -{ 1'b0,x56 } )+$signed( { 2'b0,x57 } <<<3'd1 )+$signed( { 3'b0,x58 }<<<3'd2 )+$signed( -{ 3'b0,x60 }<<<3'd2)+$signed( -{ 1'b0,x61 } )+$signed( { 2'b0,x62 } <<<3'd1 )+$signed( -{ 2'b0,x63 }<<<3'd1 )+$signed( { 1'b0,x64 }  )+$signed( -{ 3'b0,x65 }<<<3'd2)+$signed( -{ 3'b0,x67 }<<<3'd2)+$signed( { 3'b0,x68 }<<<3'd2 )+$signed( -{ 1'b0,x69 } )+$signed( -{ 3'b0,x70 }<<<3'd2)+$signed( -{ 3'b0,x71 }<<<3'd2)+$signed( -{ 3'b0,x72 }<<<3'd2)+$signed( { 1'b0,x74 }  )+$signed( { 2'b0,x75 } <<<3'd1 )+$signed( { 1'b0,x76 }  )+$signed( { 1'b0,x77 }  )+$signed( -{ 2'b0,x78 }<<<3'd1 )+$signed( { 2'b0,x79 } <<<3'd1 )+$signed( { 2'b0,x80 } <<<3'd1 )+$signed( -{ 2'b0,x81 }<<<3'd1 )+$signed( -{ 1'b0,x83 } )+$signed( -{ 2'b0,x84 }<<<3'd1 )+$signed( -{ 2'b0,x85 }<<<3'd1 )+$signed( -{ 1'b0,x86 } )+$signed( { 3'b0,x87 }<<<3'd2 )+$signed( { 2'b0,x88 } <<<3'd1 )+$signed( -{ 3'b0,x89 }<<<3'd2)+$signed( -{ 3'b0,x90 }<<<3'd2)+$signed( { 1'b0,x91 }  )+$signed( { 3'b0,x92 }<<<3'd2 )+$signed( { 2'b0,x93 } <<<3'd1 )+$signed( -{ 1'b0,x94 } )+$signed( -{ 2'b0,x95 }<<<3'd1 )+$signed( { 2'b0,x96 } <<<3'd1 )+$signed( -{ 2'b0,x97 }<<<3'd1 )+$signed( { 2'b0,x98 } <<<3'd1 )+$signed( { 2'b0,x99 } <<<3'd1 )+$signed( { 2'b0,x100 } <<<3'd1 )+$signed( -{ 2'b0,x101 }<<<3'd1 )+$signed( { 3'b0,x102 }<<<3'd2 )+$signed( { 1'b0,x103 }  )+$signed( -{ 1'b0,x104 } )+$signed( -{ 1'b0,x105 } )+$signed( { 1'b0,x106 }  )+$signed( { 1'b0,x107 }  )+$signed( { 2'b0,x108 } <<<3'd1 )+$signed( -{ 1'b0,x109 } )+$signed( { 2'b0,x110 } <<<3'd1 )+$signed( { 3'b0,x111 }<<<3'd2 )+$signed( { 2'b0,x112 } <<<3'd1 )+$signed( -{ 4'b0, x113 }<<<3'd3 )+$signed( { 2'b0,x114 } <<<3'd1 )+$signed( -{ 1'b0,x115 } )+$signed( { 3'b0,x116 }<<<3'd2 )+$signed( -{ 3'b0,x118 }<<<3'd2)+$signed( -{ 3'b0,x119 }<<<3'd2)+$signed( -{ 2'b0,x122 }<<<3'd1 )+$signed( -{ 2'b0,x123 }<<<3'd1 )+$signed( { 3'b0,x124 }<<<3'd2 )+$signed( { 2'b0,x125 } <<<3'd1 )+$signed( { 3'b0,x126 }<<<3'd2 )+$signed( { 1'b0,x128 }  )+$signed( -{ 2'b0,x129 }<<<3'd1 )+$signed( { 2'b0,x130 } <<<3'd1 )+$signed( { 1'b0,x131 }  )+$signed( -{ 2'b0,x132 }<<<3'd1 )+$signed( { 2'b0,x133 } <<<3'd1 )+$signed( { 3'b0,x135 }<<<3'd2 )+$signed( { 1'b0,x136 }  )+$signed( -{ 3'b0,x137 }<<<3'd2)+$signed( -{ 2'b0,x138 }<<<3'd1 )+$signed( -{ 1'b0,x139 } )+$signed( -{ 2'b0,x140 }<<<3'd1 )+$signed( { 3'b0,x142 }<<<3'd2 )+$signed( { 1'b0,x143 }  )+$signed( { 4'b0,x144 }<<<3'd3 )+$signed( -{ 3'b0,x145 }<<<3'd2)+$signed( { 2'b0,x146 } <<<3'd1 )+$signed( { 1'b0,x147 }  )+$signed( -{ 1'b0,x148 } )+$signed( -{ 3'b0,x149 }<<<3'd2)+$signed( -{ 1'b0,x151 } )+$signed( { 2'b0,x152 } <<<3'd1 )+$signed( { 3'b0,x153 }<<<3'd2 )+$signed( -{ 1'b0,x154 } )+$signed( { 3'b0,x155 }<<<3'd2 )+$signed( { 2'b0,x156 } <<<3'd1 )+$signed( { 3'b0,x157 }<<<3'd2 )+$signed( -{ 3'b0,x158 }<<<3'd2)+$signed( { 2'b0,x159 } <<<3'd1 )+$signed( { 3'b0,x160 }<<<3'd2 )+$signed( -{ 1'b0,x161 } )+$signed( { 3'b0,x163 }<<<3'd2 )+$signed( -{ 2'b0,x164 }<<<3'd1 )+$signed( { 3'b0,x165 }<<<3'd2 )+$signed( { 2'b0,x166 } <<<3'd1 )+$signed( -{ 3'b0,x167 }<<<3'd2)+$signed( -{ 4'b0, x168 }<<<3'd3 )+$signed( -{ 3'b0,x169 }<<<3'd2)+$signed( -{ 1'b0,x170 } )+$signed( { 3'b0,x171 }<<<3'd2 )+$signed( { 3'b0,x172 }<<<3'd2 )+$signed( { 2'b0,x173 } <<<3'd1 )+$signed( { 2'b0,x175 } <<<3'd1 )+$signed( { 1'b0,x176 }  )+$signed( -{ 1'b0,x177 } )+$signed( -{ 1'b0,x178 } )+$signed( { 3'b0,x180 }<<<3'd2 )+$signed( { 2'b0,x181 } <<<3'd1 )+$signed( -{ 4'b0, x183 }<<<3'd3 )+$signed( { 1'b0,x184 }  )+$signed( { 3'b0,x185 }<<<3'd2 )+$signed( -{ 4'b0, x186 }<<<3'd3 )+$signed( -{ 3'b0,x187 }<<<3'd2)+$signed( -{ 2'b0,x188 }<<<3'd1 )+$signed( { 4'b0,x189 }<<<3'd3 )+$signed( { 2'b0,x190 } <<<3'd1 )+$signed( -{ 2'b0,x192 }<<<3'd1 )+$signed( { 2'b0,x193 } <<<3'd1 )+$signed( { 2'b0,x194 } <<<3'd1 )+$signed( -{ 2'b0,x195 }<<<3'd1 )+$signed( { 1'b0,x196 }  )+$signed( -{ 2'b0,x197 }<<<3'd1 )+$signed( -{ 3'b0,x198 }<<<3'd2)+$signed( { 2'b0,x199 } <<<3'd1 )+$signed( -{ 2'b0,x200 }<<<3'd1 )+$signed( { 3'b0,x201 }<<<3'd2 )+$signed( { 3'b0,x202 }<<<3'd2 )+$signed( -{ 3'b0,x203 }<<<3'd2)+$signed( -{ 4'b0, x204 }<<<3'd3 )+$signed( { 3'b0,x205 }<<<3'd2 )+$signed( -{ 3'b0,x206 }<<<3'd2)+$signed( { 2'b0,x207 } <<<3'd1 )+$signed( -{ 2'b0,x208 }<<<3'd1 )+$signed( -{ 1'b0,x209 } )+$signed( { 1'b0,x210 }  )+$signed( -{ 2'b0,x211 }<<<3'd1 )+$signed( { 3'b0,x212 }<<<3'd2 )+$signed( -{ 3'b0,x213 }<<<3'd2)+$signed( -{ 3'b0,x214 }<<<3'd2)+$signed( { 3'b0,x215 }<<<3'd2 )+$signed( { 2'b0,x216 } <<<3'd1 )+$signed( { 2'b0,x217 } <<<3'd1 )+$signed( -{ 3'b0,x218 }<<<3'd2)+$signed( { 3'b0,x219 }<<<3'd2 )+$signed( { 3'b0,x220 }<<<3'd2 )+$signed( -{ 1'b0,x221 } )+$signed( -{ 3'b0,x222 }<<<3'd2)+$signed( -{ 2'b0,x223 }<<<3'd1 )+$signed( -{ 3'b0,x226 }<<<3'd2)+$signed( -{ 1'b0,x227 } )+$signed( -{ 3'b0,x228 }<<<3'd2)+$signed( -{ 3'b0,x230 }<<<3'd2)+$signed( { 1'b0,x231 }  )+$signed( -{ 3'b0,x232 }<<<3'd2)+$signed( { 2'b0,x233 } <<<3'd1 )+$signed( -{ 1'b0,x234 } )+$signed( { 3'b0,x235 }<<<3'd2 )+$signed( { 3'b0,x236 }<<<3'd2 )+$signed( { 3'b0,x237 }<<<3'd2 )+$signed( { 3'b0,x238 }<<<3'd2 )+$signed( { 1'b0,x239 }  )+$signed( -{ 4'b0, x240 }<<<3'd3 )+$signed( { 3'b0,x241 }<<<3'd2 )+$signed( -{ 3'b0,x242 }<<<3'd2)+$signed( -{ 3'b0,x243 }<<<3'd2)+$signed( -{ 2'b0,x244 }<<<3'd1 )+$signed( { 1'b0,x245 }  )+$signed( -{ 1'b0,x246 } )+$signed( -{ 4'b0, x247 }<<<3'd3 )+$signed( { 1'b0,x248 }  )+$signed( -{ 2'b0,x249 }<<<3'd1 )+$signed( { 2'b0,x251 } <<<3'd1 )+$signed( -{ 1'b0,x252 } )+$signed( { 1'b0,x253 }  )+$signed( -{ 3'b0,x254 }<<<3'd2)+$signed( -{ 1'b0,x255 } )+$signed( -{ 3'b0,x256 }<<<3'd2)+$signed( { 2'b0,x257 } <<<3'd1 )+$signed( -{ 5'b0,x258 }<<<3'd4 )+$signed( { 2'b0,x259 } <<<3'd1 )+$signed( -{ 3'b0,x260 }<<<3'd2)+$signed( { 2'b0,x261 } <<<3'd1 )+$signed( -{ 3'b0,x263 }<<<3'd2)+$signed( -{ 3'b0,x264 }<<<3'd2)+$signed( -{ 3'b0,x266 }<<<3'd2)+$signed( { 1'b0,x267 }  )+$signed( { 2'b0,x268 } <<<3'd1 )+$signed( { 2'b0,x269 } <<<3'd1 )+$signed( -{ 2'b0,x270 }<<<3'd1 )+$signed( { 3'b0,x271 }<<<3'd2 )+$signed( { 1'b0,x272 }  )+$signed( -{ 2'b0,x273 }<<<3'd1 )+$signed( { 3'b0,x274 }<<<3'd2 )+$signed( -{ 3'b0,x275 }<<<3'd2)+$signed( -{ 3'b0,x276 }<<<3'd2)+$signed( { 2'b0,x277 } <<<3'd1 )+$signed( -{ 1'b0,x278 } )+$signed( -{ 2'b0,x279 }<<<3'd1 )+$signed( -{ 3'b0,x280 }<<<3'd2)+$signed( { 2'b0,x281 } <<<3'd1 )+$signed( { 3'b0,x282 }<<<3'd2 )+$signed( -{ 4'b0, x284 }<<<3'd3 )+$signed( -{ 4'b0, x285 }<<<3'd3 )+$signed( { 2'b0,x286 } <<<3'd1 )+$signed( { 3'b0,x287 }<<<3'd2 )+$signed( { 3'b0,x289 }<<<3'd2 )+$signed( -{ 4'b0, x291 }<<<3'd3 )+$signed( { 2'b0,x292 } <<<3'd1 )+$signed( { 2'b0,x293 } <<<3'd1 )+$signed( -{ 3'b0,x294 }<<<3'd2)+$signed( -{ 3'b0,x295 }<<<3'd2)+$signed( { 1'b0,x296 }  )+$signed( { 2'b0,x299 } <<<3'd1 )+$signed( { 3'b0,x300 }<<<3'd2 )+$signed( { 2'b0,x301 } <<<3'd1 )+$signed( { 2'b0,x302 } <<<3'd1 )+$signed( -{ 2'b0,x303 }<<<3'd1 )+$signed( -{ 4'b0, x304 }<<<3'd3 )+$signed( { 3'b0,x305 }<<<3'd2 )+$signed( -{ 1'b0,x306 } )+$signed( { 2'b0,x307 } <<<3'd1 )+$signed( -{ 4'b0, x308 }<<<3'd3 )+$signed( -{ 2'b0,x309 }<<<3'd1 )+$signed( { 3'b0,x311 }<<<3'd2 )+$signed( { 3'b0,x312 }<<<3'd2 )+$signed( { 3'b0,x313 }<<<3'd2 )+$signed( { 4'b0,x314 }<<<3'd3 )+$signed( -{ 3'b0,x315 }<<<3'd2)+$signed( -{ 4'b0, x317 }<<<3'd3 )+$signed( -{ 2'b0,x318 }<<<3'd1 )+$signed( { 1'b0,x319 }  )+$signed( { 1'b0,x320 }  )+$signed( -{ 4'b0, x321 }<<<3'd3 )+$signed( { 1'b0,x323 }  )+$signed( { 3'b0,x325 }<<<3'd2 )+$signed( { 3'b0,x326 }<<<3'd2 )+$signed( -{ 3'b0,x327 }<<<3'd2)+$signed( -{ 1'b0,x328 } )+$signed( { 2'b0,x329 } <<<3'd1 )+$signed( -{ 4'b0, x330 }<<<3'd3 )+$signed( { 3'b0,x331 }<<<3'd2 )+$signed( -{ 1'b0,x332 } )+$signed( { 3'b0,x333 }<<<3'd2 )+$signed( -{ 3'b0,x334 }<<<3'd2)+$signed( { 3'b0,x335 }<<<3'd2 )+$signed( -{ 3'b0,x336 }<<<3'd2)+$signed( { 2'b0,x337 } <<<3'd1 )+$signed( -{ 3'b0,x338 }<<<3'd2)+$signed( { 3'b0,x339 }<<<3'd2 )+$signed( -{ 2'b0,x340 }<<<3'd1 )+$signed( { 2'b0,x341 } <<<3'd1 )+$signed( { 3'b0,x342 }<<<3'd2 )+$signed( -{ 3'b0,x343 }<<<3'd2)+$signed( -{ 3'b0,x344 }<<<3'd2)+$signed( { 3'b0,x345 }<<<3'd2 )+$signed( -{ 3'b0,x347 }<<<3'd2)+$signed( -{ 3'b0,x348 }<<<3'd2)+$signed( { 2'b0,x349 } <<<3'd1 )+$signed( { 3'b0,x350 }<<<3'd2 )+$signed( { 4'b0,x351 }<<<3'd3 )+$signed( { 2'b0,x352 } <<<3'd1 )+$signed( -{ 3'b0,x353 }<<<3'd2)+$signed( { 3'b0,x355 }<<<3'd2 )+$signed( -{ 3'b0,x356 }<<<3'd2)+$signed( { 3'b0,x357 }<<<3'd2 )+$signed( -{ 3'b0,x358 }<<<3'd2)+$signed( { 2'b0,x359 } <<<3'd1 )+$signed( -{ 1'b0,x360 } )+$signed( -{ 1'b0,x361 } )+$signed( -{ 1'b0,x363 } )+$signed( { 4'b0,x364 }<<<3'd3 )+$signed( -{ 3'b0,x365 }<<<3'd2)+$signed( -{ 3'b0,x366 }<<<3'd2)+$signed( -{ 2'b0,x367 }<<<3'd1 )+$signed( -{ 3'b0,x368 }<<<3'd2)+$signed( -{ 4'b0, x369 }<<<3'd3 )+$signed( { 3'b0,x370 }<<<3'd2 )+$signed( { 3'b0,x371 }<<<3'd2 )+$signed( { 1'b0,x373 }  )+$signed( -{ 1'b0,x374 } )+$signed( { 3'b0,x375 }<<<3'd2 )+$signed( -{ 1'b0,x376 } )+$signed( { 1'b0,x377 }  )+$signed( -{ 4'b0, x379 }<<<3'd3 )+$signed( -{ 3'b0,x380 }<<<3'd2)+$signed( -{ 2'b0,x381 }<<<3'd1 )+$signed( -{ 2'b0,x382 }<<<3'd1 )+$signed( -{ 2'b0,x383 }<<<3'd1 )+$signed( { 2'b0,x384 } <<<3'd1 )+$signed( { 3'b0,x385 }<<<3'd2 )+$signed( -{ 3'b0,x386 }<<<3'd2)+$signed( { 3'b0,x387 }<<<3'd2 )+$signed( { 2'b0,x388 } <<<3'd1 )+$signed( { 3'b0,x389 }<<<3'd2 )+$signed( -{ 3'b0,x390 }<<<3'd2)+$signed( { 3'b0,x391 }<<<3'd2 )+$signed( -{ 2'b0,x393 }<<<3'd1 )+$signed( -{ 1'b0,x394 } )+$signed( -{ 3'b0,x395 }<<<3'd2)+$signed( -{ 4'b0, x396 }<<<3'd3 )+$signed( { 3'b0,x397 }<<<3'd2 )+$signed( -{ 2'b0,x398 }<<<3'd1 )+$signed( -{ 2'b0,x399 }<<<3'd1 )+$signed( -{ 3'b0,x400 }<<<3'd2)+$signed( -{ 1'b0,x401 } )+$signed( { 2'b0,x402 } <<<3'd1 )+$signed( { 1'b0,x404 }  )+$signed( -{ 1'b0,x405 } )+$signed( { 3'b0,x406 }<<<3'd2 )+$signed( -{ 4'b0, x407 }<<<3'd3 )+$signed( -{ 1'b0,x408 } )+$signed( { 3'b0,x410 }<<<3'd2 )+$signed( -{ 2'b0,x411 }<<<3'd1 )+$signed( { 1'b0,x412 }  )+$signed( -{ 5'b0,x413 }<<<3'd4 )+$signed( { 3'b0,x414 }<<<3'd2 )+$signed( -{ 4'b0, x415 }<<<3'd3 )+$signed( -{ 4'b0, x416 }<<<3'd3 )+$signed( { 1'b0,x417 }  )+$signed( { 2'b0,x418 } <<<3'd1 )+$signed( { 3'b0,x419 }<<<3'd2 )+$signed( -{ 3'b0,x420 }<<<3'd2)+$signed( { 3'b0,x421 }<<<3'd2 )+$signed( { 2'b0,x422 } <<<3'd1 )+$signed( { 2'b0,x423 } <<<3'd1 )+$signed( { 3'b0,x425 }<<<3'd2 )+$signed( { 2'b0,x426 } <<<3'd1 )+$signed( -{ 4'b0, x427 }<<<3'd3 )+$signed( -{ 1'b0,x428 } )+$signed( -{ 3'b0,x429 }<<<3'd2)+$signed( -{ 2'b0,x430 }<<<3'd1 )+$signed( -{ 3'b0,x431 }<<<3'd2)+$signed( { 2'b0,x433 } <<<3'd1 )+$signed( { 2'b0,x435 } <<<3'd1 )+$signed( -{ 3'b0,x436 }<<<3'd2)+$signed( -{ 1'b0,x437 } )+$signed( -{ 4'b0, x438 }<<<3'd3 )+$signed( { 3'b0,x439 }<<<3'd2 )+$signed( { 1'b0,x440 }  )+$signed( { 1'b0,x441 }  )+$signed( { 1'b0,x442 }  )+$signed( { 3'b0,x443 }<<<3'd2 )+$signed( { 2'b0,x446 } <<<3'd1 )+$signed( -{ 3'b0,x447 }<<<3'd2)+$signed( { 3'b0,x448 }<<<3'd2 )+$signed( { 2'b0,x449 } <<<3'd1 )+$signed( { 2'b0,x450 } <<<3'd1 )+$signed( -{ 3'b0,x451 }<<<3'd2)+$signed( { 2'b0,x452 } <<<3'd1 )+$signed( -{ 1'b0,x453 } )+$signed( -{ 4'b0, x455 }<<<3'd3 )+$signed( { 1'b0,x456 }  )+$signed( { 3'b0,x457 }<<<3'd2 )+$signed( -{ 4'b0, x458 }<<<3'd3 )+$signed( { 2'b0,x459 } <<<3'd1 )+$signed( -{ 4'b0, x460 }<<<3'd3 )+$signed( -{ 2'b0,x461 }<<<3'd1 )+$signed( { 1'b0,x462 }  )+$signed( -{ 2'b0,x463 }<<<3'd1 )+$signed( -{ 2'b0,x464 }<<<3'd1 )+$signed( -{ 2'b0,x465 }<<<3'd1 )+$signed( -{ 3'b0,x466 }<<<3'd2)+$signed( -{ 4'b0, x467 }<<<3'd3 )+$signed( -{ 4'b0, x468 }<<<3'd3 )+$signed( { 3'b0,x469 }<<<3'd2 )+$signed( -{ 1'b0,x470 } )+$signed( -{ 4'b0, x471 }<<<3'd3 )+$signed( { 3'b0,x472 }<<<3'd2 )+$signed( -{ 3'b0,x473 }<<<3'd2)+$signed( -{ 3'b0,x474 }<<<3'd2)+$signed( { 3'b0,x475 }<<<3'd2 )+$signed( -{ 3'b0,x476 }<<<3'd2)+$signed( { 3'b0,x477 }<<<3'd2 )+$signed( -{ 4'b0, x478 }<<<3'd3 )+$signed( -{ 2'b0,x480 }<<<3'd1 )+$signed( -{ 3'b0,x481 }<<<3'd2)+$signed( { 2'b0,x482 } <<<3'd1 )+$signed( { 2'b0,x484 } <<<3'd1 )+$signed( { 2'b0,x485 } <<<3'd1 )+$signed( -{ 3'b0,x486 }<<<3'd2)+$signed( { 3'b0,x487 }<<<3'd2 )+$signed( { 2'b0,x488 } <<<3'd1 )+$signed( { 1'b0,x489 }  )+$signed( -{ 3'b0,x490 }<<<3'd2)+$signed( -{ 2'b0,x491 }<<<3'd1 )+$signed( -{ 3'b0,x492 }<<<3'd2)+$signed( { 2'b0,x493 } <<<3'd1 )+$signed( -{ 2'b0,x494 }<<<3'd1 )+$signed( { 4'b0,x495 }<<<3'd3 )-$signed(13'd8);
assign y17=temp_y[17][13] ==1'b1 ? 6'd0 :  
    temp_y[17][10] ==1'b1 ? 6'd63 : 
    temp_y[17][3]==1'b1 ? temp_y[17][9:4]+1'b1 : temp_y[17][9:4];
assign temp_y[18] = 
+$signed( -{ 3'b0,x0 }<<<3'd2)+$signed( -{ 3'b0,x2 }<<<3'd2)+$signed( { 3'b0,x3 }<<<3'd2 )+$signed( -{ 1'b0,x4 } )+$signed( -{ 1'b0,x5 } )+$signed( { 2'b0,x7 } <<<3'd1 )+$signed( -{ 2'b0,x9 }<<<3'd1 )+$signed( { 3'b0,x12 }<<<3'd2 )+$signed( { 1'b0,x13 }  )+$signed( { 2'b0,x14 } <<<3'd1 )+$signed( { 1'b0,x15 }  )+$signed( -{ 3'b0,x16 }<<<3'd2)+$signed( -{ 1'b0,x17 } )+$signed( -{ 3'b0,x18 }<<<3'd2)+$signed( -{ 1'b0,x19 } )+$signed( -{ 2'b0,x20 }<<<3'd1 )+$signed( -{ 1'b0,x21 } )+$signed( -{ 1'b0,x22 } )+$signed( -{ 2'b0,x23 }<<<3'd1 )+$signed( -{ 3'b0,x24 }<<<3'd2)+$signed( -{ 1'b0,x25 } )+$signed( { 2'b0,x26 } <<<3'd1 )+$signed( -{ 3'b0,x27 }<<<3'd2)+$signed( { 4'b0,x28 }<<<3'd3 )+$signed( -{ 2'b0,x30 }<<<3'd1 )+$signed( -{ 1'b0,x31 } )+$signed( -{ 1'b0,x32 } )+$signed( { 1'b0,x33 }  )+$signed( -{ 3'b0,x34 }<<<3'd2)+$signed( -{ 1'b0,x35 } )+$signed( { 2'b0,x36 } <<<3'd1 )+$signed( { 2'b0,x37 } <<<3'd1 )+$signed( -{ 3'b0,x38 }<<<3'd2)+$signed( -{ 3'b0,x39 }<<<3'd2)+$signed( -{ 1'b0,x40 } )+$signed( -{ 4'b0, x41 }<<<3'd3 )+$signed( -{ 2'b0,x42 }<<<3'd1 )+$signed( { 2'b0,x43 } <<<3'd1 )+$signed( { 2'b0,x45 } <<<3'd1 )+$signed( { 2'b0,x46 } <<<3'd1 )+$signed( -{ 1'b0,x47 } )+$signed( -{ 2'b0,x48 }<<<3'd1 )+$signed( -{ 1'b0,x50 } )+$signed( -{ 1'b0,x51 } )+$signed( -{ 1'b0,x52 } )+$signed( { 1'b0,x53 }  )+$signed( -{ 1'b0,x55 } )+$signed( { 2'b0,x56 } <<<3'd1 )+$signed( -{ 2'b0,x58 }<<<3'd1 )+$signed( { 2'b0,x59 } <<<3'd1 )+$signed( { 2'b0,x60 } <<<3'd1 )+$signed( -{ 2'b0,x62 }<<<3'd1 )+$signed( -{ 2'b0,x63 }<<<3'd1 )+$signed( -{ 2'b0,x64 }<<<3'd1 )+$signed( -{ 2'b0,x66 }<<<3'd1 )+$signed( { 3'b0,x67 }<<<3'd2 )+$signed( { 2'b0,x68 } <<<3'd1 )+$signed( { 3'b0,x69 }<<<3'd2 )+$signed( -{ 2'b0,x70 }<<<3'd1 )+$signed( -{ 4'b0, x71 }<<<3'd3 )+$signed( -{ 2'b0,x72 }<<<3'd1 )+$signed( -{ 2'b0,x75 }<<<3'd1 )+$signed( { 2'b0,x76 } <<<3'd1 )+$signed( { 2'b0,x77 } <<<3'd1 )+$signed( -{ 1'b0,x78 } )+$signed( -{ 3'b0,x80 }<<<3'd2)+$signed( { 3'b0,x81 }<<<3'd2 )+$signed( -{ 3'b0,x82 }<<<3'd2)+$signed( -{ 3'b0,x83 }<<<3'd2)+$signed( { 3'b0,x84 }<<<3'd2 )+$signed( { 1'b0,x85 }  )+$signed( { 3'b0,x87 }<<<3'd2 )+$signed( { 2'b0,x88 } <<<3'd1 )+$signed( -{ 2'b0,x89 }<<<3'd1 )+$signed( { 4'b0,x90 }<<<3'd3 )+$signed( -{ 2'b0,x91 }<<<3'd1 )+$signed( { 3'b0,x93 }<<<3'd2 )+$signed( -{ 3'b0,x94 }<<<3'd2)+$signed( { 2'b0,x96 } <<<3'd1 )+$signed( -{ 4'b0, x97 }<<<3'd3 )+$signed( { 3'b0,x98 }<<<3'd2 )+$signed( -{ 1'b0,x100 } )+$signed( -{ 1'b0,x101 } )+$signed( { 3'b0,x102 }<<<3'd2 )+$signed( { 3'b0,x103 }<<<3'd2 )+$signed( { 3'b0,x104 }<<<3'd2 )+$signed( -{ 2'b0,x105 }<<<3'd1 )+$signed( -{ 3'b0,x106 }<<<3'd2)+$signed( { 3'b0,x107 }<<<3'd2 )+$signed( { 1'b0,x108 }  )+$signed( -{ 2'b0,x109 }<<<3'd1 )+$signed( { 1'b0,x110 }  )+$signed( -{ 1'b0,x111 } )+$signed( { 2'b0,x112 } <<<3'd1 )+$signed( { 4'b0,x115 }<<<3'd3 )+$signed( -{ 3'b0,x116 }<<<3'd2)+$signed( -{ 3'b0,x117 }<<<3'd2)+$signed( { 2'b0,x118 } <<<3'd1 )+$signed( { 3'b0,x119 }<<<3'd2 )+$signed( -{ 4'b0, x120 }<<<3'd3 )+$signed( -{ 3'b0,x121 }<<<3'd2)+$signed( { 2'b0,x122 } <<<3'd1 )+$signed( -{ 3'b0,x123 }<<<3'd2)+$signed( -{ 1'b0,x124 } )+$signed( { 1'b0,x126 }  )+$signed( -{ 3'b0,x127 }<<<3'd2)+$signed( -{ 1'b0,x128 } )+$signed( -{ 1'b0,x130 } )+$signed( { 1'b0,x131 }  )+$signed( -{ 3'b0,x133 }<<<3'd2)+$signed( -{ 1'b0,x134 } )+$signed( { 2'b0,x135 } <<<3'd1 )+$signed( { 3'b0,x136 }<<<3'd2 )+$signed( { 2'b0,x138 } <<<3'd1 )+$signed( -{ 3'b0,x139 }<<<3'd2)+$signed( -{ 1'b0,x140 } )+$signed( { 3'b0,x141 }<<<3'd2 )+$signed( { 3'b0,x142 }<<<3'd2 )+$signed( -{ 4'b0, x143 }<<<3'd3 )+$signed( { 1'b0,x144 }  )+$signed( -{ 3'b0,x145 }<<<3'd2)+$signed( { 3'b0,x146 }<<<3'd2 )+$signed( -{ 3'b0,x147 }<<<3'd2)+$signed( -{ 2'b0,x148 }<<<3'd1 )+$signed( -{ 1'b0,x149 } )+$signed( -{ 3'b0,x150 }<<<3'd2)+$signed( { 2'b0,x151 } <<<3'd1 )+$signed( -{ 3'b0,x152 }<<<3'd2)+$signed( { 2'b0,x153 } <<<3'd1 )+$signed( -{ 3'b0,x154 }<<<3'd2)+$signed( -{ 3'b0,x155 }<<<3'd2)+$signed( -{ 4'b0, x156 }<<<3'd3 )+$signed( -{ 3'b0,x157 }<<<3'd2)+$signed( { 2'b0,x158 } <<<3'd1 )+$signed( { 3'b0,x159 }<<<3'd2 )+$signed( -{ 2'b0,x160 }<<<3'd1 )+$signed( -{ 3'b0,x161 }<<<3'd2)+$signed( { 3'b0,x162 }<<<3'd2 )+$signed( -{ 3'b0,x163 }<<<3'd2)+$signed( -{ 2'b0,x164 }<<<3'd1 )+$signed( -{ 1'b0,x165 } )+$signed( -{ 4'b0, x166 }<<<3'd3 )+$signed( { 2'b0,x169 } <<<3'd1 )+$signed( { 2'b0,x170 } <<<3'd1 )+$signed( -{ 3'b0,x171 }<<<3'd2)+$signed( -{ 1'b0,x173 } )+$signed( { 2'b0,x174 } <<<3'd1 )+$signed( { 4'b0,x176 }<<<3'd3 )+$signed( { 3'b0,x177 }<<<3'd2 )+$signed( -{ 1'b0,x178 } )+$signed( -{ 2'b0,x179 }<<<3'd1 )+$signed( -{ 1'b0,x180 } )+$signed( -{ 4'b0, x181 }<<<3'd3 )+$signed( { 4'b0,x182 }<<<3'd3 )+$signed( { 3'b0,x183 }<<<3'd2 )+$signed( { 3'b0,x184 }<<<3'd2 )+$signed( { 1'b0,x185 }  )+$signed( { 3'b0,x186 }<<<3'd2 )+$signed( { 2'b0,x187 } <<<3'd1 )+$signed( -{ 2'b0,x188 }<<<3'd1 )+$signed( -{ 4'b0, x190 }<<<3'd3 )+$signed( -{ 3'b0,x191 }<<<3'd2)+$signed( -{ 3'b0,x193 }<<<3'd2)+$signed( -{ 3'b0,x194 }<<<3'd2)+$signed( { 3'b0,x195 }<<<3'd2 )+$signed( -{ 3'b0,x196 }<<<3'd2)+$signed( -{ 4'b0, x197 }<<<3'd3 )+$signed( -{ 3'b0,x198 }<<<3'd2)+$signed( -{ 2'b0,x199 }<<<3'd1 )+$signed( -{ 3'b0,x200 }<<<3'd2)+$signed( { 3'b0,x201 }<<<3'd2 )+$signed( -{ 3'b0,x202 }<<<3'd2)+$signed( -{ 4'b0, x203 }<<<3'd3 )+$signed( { 2'b0,x204 } <<<3'd1 )+$signed( -{ 4'b0, x205 }<<<3'd3 )+$signed( { 3'b0,x206 }<<<3'd2 )+$signed( -{ 3'b0,x207 }<<<3'd2)+$signed( { 4'b0,x208 }<<<3'd3 )+$signed( -{ 1'b0,x209 } )+$signed( { 1'b0,x210 }  )+$signed( -{ 1'b0,x211 } )+$signed( { 4'b0,x212 }<<<3'd3 )+$signed( -{ 1'b0,x213 } )+$signed( { 3'b0,x214 }<<<3'd2 )+$signed( { 3'b0,x215 }<<<3'd2 )+$signed( { 2'b0,x216 } <<<3'd1 )+$signed( -{ 4'b0, x217 }<<<3'd3 )+$signed( { 3'b0,x218 }<<<3'd2 )+$signed( -{ 3'b0,x220 }<<<3'd2)+$signed( { 2'b0,x221 } <<<3'd1 )+$signed( { 3'b0,x222 }<<<3'd2 )+$signed( -{ 3'b0,x223 }<<<3'd2)+$signed( { 1'b0,x224 }  )+$signed( -{ 3'b0,x225 }<<<3'd2)+$signed( -{ 1'b0,x226 } )+$signed( { 2'b0,x227 } <<<3'd1 )+$signed( -{ 2'b0,x228 }<<<3'd1 )+$signed( -{ 1'b0,x230 } )+$signed( { 3'b0,x231 }<<<3'd2 )+$signed( -{ 4'b0, x232 }<<<3'd3 )+$signed( -{ 1'b0,x233 } )+$signed( -{ 3'b0,x234 }<<<3'd2)+$signed( { 2'b0,x235 } <<<3'd1 )+$signed( -{ 3'b0,x236 }<<<3'd2)+$signed( { 3'b0,x237 }<<<3'd2 )+$signed( -{ 3'b0,x238 }<<<3'd2)+$signed( { 2'b0,x239 } <<<3'd1 )+$signed( { 1'b0,x240 }  )+$signed( -{ 4'b0, x241 }<<<3'd3 )+$signed( { 2'b0,x242 } <<<3'd1 )+$signed( -{ 2'b0,x243 }<<<3'd1 )+$signed( { 2'b0,x244 } <<<3'd1 )+$signed( { 2'b0,x245 } <<<3'd1 )+$signed( -{ 3'b0,x246 }<<<3'd2)+$signed( { 3'b0,x248 }<<<3'd2 )+$signed( -{ 3'b0,x250 }<<<3'd2)+$signed( { 3'b0,x251 }<<<3'd2 )+$signed( -{ 1'b0,x252 } )+$signed( -{ 3'b0,x253 }<<<3'd2)+$signed( { 3'b0,x254 }<<<3'd2 )+$signed( -{ 1'b0,x255 } )+$signed( { 1'b0,x256 }  )+$signed( -{ 1'b0,x257 } )+$signed( { 2'b0,x258 } <<<3'd1 )+$signed( -{ 2'b0,x259 }<<<3'd1 )+$signed( -{ 2'b0,x260 }<<<3'd1 )+$signed( -{ 1'b0,x261 } )+$signed( -{ 1'b0,x262 } )+$signed( { 1'b0,x263 }  )+$signed( -{ 3'b0,x264 }<<<3'd2)+$signed( { 1'b0,x265 }  )+$signed( { 1'b0,x266 }  )+$signed( { 2'b0,x267 } <<<3'd1 )+$signed( -{ 2'b0,x268 }<<<3'd1 )+$signed( { 3'b0,x270 }<<<3'd2 )+$signed( { 2'b0,x271 } <<<3'd1 )+$signed( -{ 3'b0,x272 }<<<3'd2)+$signed( { 4'b0,x273 }<<<3'd3 )+$signed( -{ 3'b0,x274 }<<<3'd2)+$signed( -{ 4'b0, x277 }<<<3'd3 )+$signed( { 3'b0,x278 }<<<3'd2 )+$signed( -{ 3'b0,x279 }<<<3'd2)+$signed( -{ 3'b0,x280 }<<<3'd2)+$signed( -{ 2'b0,x281 }<<<3'd1 )+$signed( { 1'b0,x283 }  )+$signed( { 4'b0,x284 }<<<3'd3 )+$signed( -{ 3'b0,x285 }<<<3'd2)+$signed( -{ 1'b0,x286 } )+$signed( { 3'b0,x287 }<<<3'd2 )+$signed( { 3'b0,x289 }<<<3'd2 )+$signed( -{ 1'b0,x290 } )+$signed( { 2'b0,x291 } <<<3'd1 )+$signed( -{ 3'b0,x292 }<<<3'd2)+$signed( { 2'b0,x293 } <<<3'd1 )+$signed( -{ 2'b0,x294 }<<<3'd1 )+$signed( -{ 3'b0,x298 }<<<3'd2)+$signed( -{ 3'b0,x299 }<<<3'd2)+$signed( { 2'b0,x300 } <<<3'd1 )+$signed( -{ 2'b0,x301 }<<<3'd1 )+$signed( -{ 3'b0,x302 }<<<3'd2)+$signed( -{ 1'b0,x304 } )+$signed( -{ 3'b0,x305 }<<<3'd2)+$signed( { 1'b0,x306 }  )+$signed( -{ 2'b0,x307 }<<<3'd1 )+$signed( -{ 1'b0,x308 } )+$signed( -{ 4'b0, x309 }<<<3'd3 )+$signed( { 2'b0,x310 } <<<3'd1 )+$signed( { 3'b0,x311 }<<<3'd2 )+$signed( -{ 1'b0,x312 } )+$signed( { 3'b0,x313 }<<<3'd2 )+$signed( -{ 1'b0,x314 } )+$signed( -{ 2'b0,x317 }<<<3'd1 )+$signed( -{ 2'b0,x318 }<<<3'd1 )+$signed( -{ 1'b0,x319 } )+$signed( { 1'b0,x320 }  )+$signed( { 3'b0,x321 }<<<3'd2 )+$signed( { 3'b0,x322 }<<<3'd2 )+$signed( -{ 2'b0,x323 }<<<3'd1 )+$signed( -{ 3'b0,x324 }<<<3'd2)+$signed( -{ 2'b0,x325 }<<<3'd1 )+$signed( -{ 1'b0,x326 } )+$signed( -{ 3'b0,x327 }<<<3'd2)+$signed( { 3'b0,x328 }<<<3'd2 )+$signed( -{ 2'b0,x329 }<<<3'd1 )+$signed( -{ 3'b0,x330 }<<<3'd2)+$signed( { 4'b0,x331 }<<<3'd3 )+$signed( -{ 2'b0,x332 }<<<3'd1 )+$signed( { 2'b0,x333 } <<<3'd1 )+$signed( { 3'b0,x334 }<<<3'd2 )+$signed( { 3'b0,x335 }<<<3'd2 )+$signed( -{ 1'b0,x336 } )+$signed( -{ 1'b0,x338 } )+$signed( -{ 3'b0,x339 }<<<3'd2)+$signed( { 3'b0,x340 }<<<3'd2 )+$signed( { 3'b0,x341 }<<<3'd2 )+$signed( { 2'b0,x342 } <<<3'd1 )+$signed( -{ 4'b0, x343 }<<<3'd3 )+$signed( { 2'b0,x344 } <<<3'd1 )+$signed( -{ 2'b0,x345 }<<<3'd1 )+$signed( { 1'b0,x346 }  )+$signed( -{ 2'b0,x347 }<<<3'd1 )+$signed( -{ 2'b0,x348 }<<<3'd1 )+$signed( -{ 3'b0,x349 }<<<3'd2)+$signed( -{ 2'b0,x350 }<<<3'd1 )+$signed( { 1'b0,x351 }  )+$signed( { 1'b0,x352 }  )+$signed( { 2'b0,x353 } <<<3'd1 )+$signed( { 3'b0,x355 }<<<3'd2 )+$signed( { 4'b0,x356 }<<<3'd3 )+$signed( { 4'b0,x357 }<<<3'd3 )+$signed( -{ 1'b0,x359 } )+$signed( -{ 2'b0,x360 }<<<3'd1 )+$signed( { 4'b0,x361 }<<<3'd3 )+$signed( { 1'b0,x362 }  )+$signed( -{ 3'b0,x363 }<<<3'd2)+$signed( { 1'b0,x364 }  )+$signed( -{ 3'b0,x365 }<<<3'd2)+$signed( -{ 3'b0,x366 }<<<3'd2)+$signed( { 2'b0,x367 } <<<3'd1 )+$signed( -{ 2'b0,x368 }<<<3'd1 )+$signed( { 2'b0,x369 } <<<3'd1 )+$signed( -{ 3'b0,x370 }<<<3'd2)+$signed( -{ 3'b0,x371 }<<<3'd2)+$signed( { 3'b0,x372 }<<<3'd2 )+$signed( { 4'b0,x375 }<<<3'd3 )+$signed( -{ 2'b0,x376 }<<<3'd1 )+$signed( -{ 4'b0, x377 }<<<3'd3 )+$signed( { 3'b0,x378 }<<<3'd2 )+$signed( { 2'b0,x379 } <<<3'd1 )+$signed( { 1'b0,x380 }  )+$signed( -{ 1'b0,x381 } )+$signed( -{ 4'b0, x383 }<<<3'd3 )+$signed( { 1'b0,x384 }  )+$signed( { 2'b0,x385 } <<<3'd1 )+$signed( { 4'b0,x386 }<<<3'd3 )+$signed( -{ 2'b0,x387 }<<<3'd1 )+$signed( -{ 1'b0,x388 } )+$signed( { 3'b0,x389 }<<<3'd2 )+$signed( { 2'b0,x390 } <<<3'd1 )+$signed( -{ 3'b0,x392 }<<<3'd2)+$signed( { 3'b0,x393 }<<<3'd2 )+$signed( { 3'b0,x394 }<<<3'd2 )+$signed( -{ 3'b0,x396 }<<<3'd2)+$signed( { 1'b0,x397 }  )+$signed( { 4'b0,x398 }<<<3'd3 )+$signed( { 3'b0,x399 }<<<3'd2 )+$signed( { 3'b0,x400 }<<<3'd2 )+$signed( -{ 3'b0,x401 }<<<3'd2)+$signed( { 2'b0,x402 } <<<3'd1 )+$signed( -{ 3'b0,x403 }<<<3'd2)+$signed( { 3'b0,x404 }<<<3'd2 )+$signed( { 3'b0,x405 }<<<3'd2 )+$signed( -{ 2'b0,x406 }<<<3'd1 )+$signed( -{ 1'b0,x407 } )+$signed( { 4'b0,x408 }<<<3'd3 )+$signed( { 1'b0,x410 }  )+$signed( -{ 3'b0,x411 }<<<3'd2)+$signed( -{ 1'b0,x412 } )+$signed( { 2'b0,x413 } <<<3'd1 )+$signed( { 4'b0,x414 }<<<3'd3 )+$signed( { 3'b0,x415 }<<<3'd2 )+$signed( -{ 3'b0,x416 }<<<3'd2)+$signed( -{ 4'b0, x417 }<<<3'd3 )+$signed( -{ 4'b0, x418 }<<<3'd3 )+$signed( { 3'b0,x419 }<<<3'd2 )+$signed( { 3'b0,x420 }<<<3'd2 )+$signed( -{ 4'b0, x421 }<<<3'd3 )+$signed( -{ 2'b0,x422 }<<<3'd1 )+$signed( -{ 3'b0,x423 }<<<3'd2)+$signed( { 2'b0,x424 } <<<3'd1 )+$signed( { 1'b0,x425 }  )+$signed( -{ 2'b0,x426 }<<<3'd1 )+$signed( -{ 3'b0,x427 }<<<3'd2)+$signed( { 3'b0,x428 }<<<3'd2 )+$signed( { 3'b0,x429 }<<<3'd2 )+$signed( -{ 3'b0,x430 }<<<3'd2)+$signed( { 3'b0,x431 }<<<3'd2 )+$signed( -{ 3'b0,x432 }<<<3'd2)+$signed( -{ 3'b0,x433 }<<<3'd2)+$signed( { 2'b0,x434 } <<<3'd1 )+$signed( -{ 5'b0,x435 }<<<3'd4 )+$signed( -{ 3'b0,x437 }<<<3'd2)+$signed( -{ 3'b0,x438 }<<<3'd2)+$signed( -{ 3'b0,x439 }<<<3'd2)+$signed( -{ 2'b0,x441 }<<<3'd1 )+$signed( { 1'b0,x442 }  )+$signed( -{ 1'b0,x443 } )+$signed( -{ 3'b0,x444 }<<<3'd2)+$signed( { 2'b0,x445 } <<<3'd1 )+$signed( { 1'b0,x447 }  )+$signed( -{ 3'b0,x448 }<<<3'd2)+$signed( { 1'b0,x449 }  )+$signed( { 3'b0,x450 }<<<3'd2 )+$signed( { 3'b0,x451 }<<<3'd2 )+$signed( -{ 2'b0,x452 }<<<3'd1 )+$signed( { 3'b0,x454 }<<<3'd2 )+$signed( -{ 4'b0, x455 }<<<3'd3 )+$signed( -{ 2'b0,x456 }<<<3'd1 )+$signed( { 1'b0,x457 }  )+$signed( -{ 1'b0,x458 } )+$signed( { 2'b0,x459 } <<<3'd1 )+$signed( { 2'b0,x460 } <<<3'd1 )+$signed( -{ 4'b0, x461 }<<<3'd3 )+$signed( { 3'b0,x462 }<<<3'd2 )+$signed( -{ 3'b0,x463 }<<<3'd2)+$signed( -{ 2'b0,x464 }<<<3'd1 )+$signed( -{ 1'b0,x465 } )+$signed( { 1'b0,x466 }  )+$signed( { 3'b0,x467 }<<<3'd2 )+$signed( { 3'b0,x468 }<<<3'd2 )+$signed( -{ 1'b0,x469 } )+$signed( { 2'b0,x470 } <<<3'd1 )+$signed( -{ 2'b0,x471 }<<<3'd1 )+$signed( -{ 3'b0,x472 }<<<3'd2)+$signed( -{ 1'b0,x473 } )+$signed( -{ 2'b0,x474 }<<<3'd1 )+$signed( { 1'b0,x476 }  )+$signed( { 1'b0,x477 }  )+$signed( { 3'b0,x478 }<<<3'd2 )+$signed( { 3'b0,x480 }<<<3'd2 )+$signed( -{ 3'b0,x481 }<<<3'd2)+$signed( -{ 2'b0,x482 }<<<3'd1 )+$signed( { 3'b0,x483 }<<<3'd2 )+$signed( -{ 4'b0, x484 }<<<3'd3 )+$signed( -{ 1'b0,x485 } )+$signed( { 1'b0,x486 }  )+$signed( -{ 3'b0,x487 }<<<3'd2)+$signed( -{ 3'b0,x489 }<<<3'd2)+$signed( -{ 2'b0,x490 }<<<3'd1 )+$signed( { 3'b0,x491 }<<<3'd2 )+$signed( { 1'b0,x492 }  )+$signed( -{ 4'b0, x493 }<<<3'd3 )+$signed( { 3'b0,x494 }<<<3'd2 )+$signed( -{ 3'b0,x495 }<<<3'd2)-$signed(13'd8);
assign y18=temp_y[18][13] ==1'b1 ? 6'd0 :  
    temp_y[18][10] ==1'b1 ? 6'd63 : 
    temp_y[18][3]==1'b1 ? temp_y[18][9:4]+1'b1 : temp_y[18][9:4];
assign temp_y[19] = 
+$signed( -{ 4'b0, x0 }<<<3'd3 )+$signed( -{ 5'b0,x1 }<<<3'd4 )+$signed( -{ 2'b0,x2 }<<<3'd1 )+$signed( -{ 2'b0,x3 }<<<3'd1 )+$signed( -{ 1'b0,x4 } )+$signed( { 2'b0,x5 } <<<3'd1 )+$signed( { 2'b0,x6 } <<<3'd1 )+$signed( { 2'b0,x7 } <<<3'd1 )+$signed( { 1'b0,x8 }  )+$signed( { 2'b0,x9 } <<<3'd1 )+$signed( { 3'b0,x10 }<<<3'd2 )+$signed( { 3'b0,x11 }<<<3'd2 )+$signed( -{ 2'b0,x12 }<<<3'd1 )+$signed( -{ 3'b0,x13 }<<<3'd2)+$signed( -{ 3'b0,x14 }<<<3'd2)+$signed( { 3'b0,x15 }<<<3'd2 )+$signed( { 1'b0,x16 }  )+$signed( -{ 3'b0,x17 }<<<3'd2)+$signed( -{ 2'b0,x18 }<<<3'd1 )+$signed( -{ 4'b0, x19 }<<<3'd3 )+$signed( -{ 2'b0,x20 }<<<3'd1 )+$signed( { 1'b0,x21 }  )+$signed( -{ 1'b0,x22 } )+$signed( -{ 1'b0,x23 } )+$signed( { 2'b0,x24 } <<<3'd1 )+$signed( { 2'b0,x25 } <<<3'd1 )+$signed( -{ 2'b0,x26 }<<<3'd1 )+$signed( -{ 3'b0,x27 }<<<3'd2)+$signed( -{ 3'b0,x30 }<<<3'd2)+$signed( -{ 2'b0,x31 }<<<3'd1 )+$signed( -{ 2'b0,x32 }<<<3'd1 )+$signed( -{ 1'b0,x33 } )+$signed( -{ 1'b0,x34 } )+$signed( -{ 1'b0,x35 } )+$signed( -{ 2'b0,x36 }<<<3'd1 )+$signed( -{ 4'b0, x37 }<<<3'd3 )+$signed( -{ 3'b0,x39 }<<<3'd2)+$signed( -{ 1'b0,x40 } )+$signed( { 1'b0,x42 }  )+$signed( -{ 1'b0,x44 } )+$signed( { 3'b0,x45 }<<<3'd2 )+$signed( { 3'b0,x47 }<<<3'd2 )+$signed( -{ 3'b0,x48 }<<<3'd2)+$signed( -{ 2'b0,x49 }<<<3'd1 )+$signed( -{ 2'b0,x50 }<<<3'd1 )+$signed( { 2'b0,x51 } <<<3'd1 )+$signed( -{ 1'b0,x52 } )+$signed( -{ 2'b0,x53 }<<<3'd1 )+$signed( -{ 1'b0,x54 } )+$signed( -{ 4'b0, x55 }<<<3'd3 )+$signed( -{ 3'b0,x56 }<<<3'd2)+$signed( -{ 3'b0,x57 }<<<3'd2)+$signed( -{ 3'b0,x58 }<<<3'd2)+$signed( -{ 1'b0,x59 } )+$signed( { 2'b0,x60 } <<<3'd1 )+$signed( { 1'b0,x61 }  )+$signed( { 1'b0,x62 }  )+$signed( { 1'b0,x63 }  )+$signed( { 2'b0,x64 } <<<3'd1 )+$signed( { 2'b0,x65 } <<<3'd1 )+$signed( { 2'b0,x66 } <<<3'd1 )+$signed( -{ 3'b0,x67 }<<<3'd2)+$signed( -{ 3'b0,x68 }<<<3'd2)+$signed( -{ 2'b0,x69 }<<<3'd1 )+$signed( { 3'b0,x70 }<<<3'd2 )+$signed( -{ 2'b0,x71 }<<<3'd1 )+$signed( -{ 2'b0,x72 }<<<3'd1 )+$signed( -{ 4'b0, x73 }<<<3'd3 )+$signed( -{ 3'b0,x75 }<<<3'd2)+$signed( { 1'b0,x76 }  )+$signed( -{ 3'b0,x77 }<<<3'd2)+$signed( { 3'b0,x78 }<<<3'd2 )+$signed( { 2'b0,x79 } <<<3'd1 )+$signed( { 2'b0,x80 } <<<3'd1 )+$signed( { 2'b0,x81 } <<<3'd1 )+$signed( { 2'b0,x83 } <<<3'd1 )+$signed( { 2'b0,x84 } <<<3'd1 )+$signed( -{ 3'b0,x86 }<<<3'd2)+$signed( { 1'b0,x87 }  )+$signed( -{ 1'b0,x88 } )+$signed( -{ 1'b0,x89 } )+$signed( -{ 1'b0,x90 } )+$signed( -{ 3'b0,x91 }<<<3'd2)+$signed( -{ 2'b0,x92 }<<<3'd1 )+$signed( -{ 3'b0,x93 }<<<3'd2)+$signed( { 1'b0,x95 }  )+$signed( { 3'b0,x96 }<<<3'd2 )+$signed( { 2'b0,x97 } <<<3'd1 )+$signed( { 1'b0,x98 }  )+$signed( -{ 2'b0,x100 }<<<3'd1 )+$signed( { 3'b0,x101 }<<<3'd2 )+$signed( -{ 1'b0,x102 } )+$signed( -{ 2'b0,x103 }<<<3'd1 )+$signed( -{ 2'b0,x104 }<<<3'd1 )+$signed( { 1'b0,x105 }  )+$signed( -{ 2'b0,x106 }<<<3'd1 )+$signed( -{ 2'b0,x107 }<<<3'd1 )+$signed( -{ 2'b0,x108 }<<<3'd1 )+$signed( -{ 4'b0, x109 }<<<3'd3 )+$signed( -{ 1'b0,x110 } )+$signed( { 2'b0,x111 } <<<3'd1 )+$signed( -{ 1'b0,x112 } )+$signed( { 2'b0,x113 } <<<3'd1 )+$signed( { 2'b0,x114 } <<<3'd1 )+$signed( -{ 3'b0,x115 }<<<3'd2)+$signed( -{ 1'b0,x116 } )+$signed( -{ 2'b0,x117 }<<<3'd1 )+$signed( { 2'b0,x118 } <<<3'd1 )+$signed( { 1'b0,x119 }  )+$signed( -{ 3'b0,x120 }<<<3'd2)+$signed( -{ 3'b0,x121 }<<<3'd2)+$signed( -{ 2'b0,x122 }<<<3'd1 )+$signed( -{ 2'b0,x123 }<<<3'd1 )+$signed( { 1'b0,x124 }  )+$signed( { 2'b0,x125 } <<<3'd1 )+$signed( -{ 3'b0,x126 }<<<3'd2)+$signed( -{ 3'b0,x127 }<<<3'd2)+$signed( { 1'b0,x128 }  )+$signed( -{ 4'b0, x129 }<<<3'd3 )+$signed( -{ 2'b0,x130 }<<<3'd1 )+$signed( -{ 1'b0,x131 } )+$signed( { 2'b0,x133 } <<<3'd1 )+$signed( -{ 1'b0,x134 } )+$signed( { 2'b0,x135 } <<<3'd1 )+$signed( -{ 1'b0,x136 } )+$signed( -{ 1'b0,x137 } )+$signed( { 2'b0,x138 } <<<3'd1 )+$signed( -{ 2'b0,x139 }<<<3'd1 )+$signed( -{ 1'b0,x140 } )+$signed( -{ 2'b0,x141 }<<<3'd1 )+$signed( { 3'b0,x142 }<<<3'd2 )+$signed( -{ 2'b0,x143 }<<<3'd1 )+$signed( -{ 2'b0,x144 }<<<3'd1 )+$signed( -{ 3'b0,x145 }<<<3'd2)+$signed( { 1'b0,x146 }  )+$signed( -{ 3'b0,x147 }<<<3'd2)+$signed( -{ 3'b0,x148 }<<<3'd2)+$signed( { 2'b0,x150 } <<<3'd1 )+$signed( { 3'b0,x151 }<<<3'd2 )+$signed( { 1'b0,x152 }  )+$signed( { 3'b0,x153 }<<<3'd2 )+$signed( -{ 2'b0,x154 }<<<3'd1 )+$signed( -{ 2'b0,x155 }<<<3'd1 )+$signed( -{ 2'b0,x157 }<<<3'd1 )+$signed( { 1'b0,x159 }  )+$signed( -{ 2'b0,x160 }<<<3'd1 )+$signed( -{ 4'b0, x161 }<<<3'd3 )+$signed( -{ 3'b0,x162 }<<<3'd2)+$signed( { 2'b0,x163 } <<<3'd1 )+$signed( { 1'b0,x164 }  )+$signed( -{ 4'b0, x165 }<<<3'd3 )+$signed( { 1'b0,x166 }  )+$signed( { 2'b0,x168 } <<<3'd1 )+$signed( { 2'b0,x169 } <<<3'd1 )+$signed( { 2'b0,x170 } <<<3'd1 )+$signed( -{ 2'b0,x171 }<<<3'd1 )+$signed( { 1'b0,x172 }  )+$signed( { 1'b0,x173 }  )+$signed( -{ 1'b0,x174 } )+$signed( { 1'b0,x175 }  )+$signed( -{ 1'b0,x176 } )+$signed( { 3'b0,x177 }<<<3'd2 )+$signed( { 2'b0,x178 } <<<3'd1 )+$signed( { 1'b0,x179 }  )+$signed( -{ 2'b0,x180 }<<<3'd1 )+$signed( { 2'b0,x181 } <<<3'd1 )+$signed( -{ 1'b0,x182 } )+$signed( { 3'b0,x183 }<<<3'd2 )+$signed( -{ 3'b0,x184 }<<<3'd2)+$signed( { 2'b0,x185 } <<<3'd1 )+$signed( { 2'b0,x186 } <<<3'd1 )+$signed( { 1'b0,x187 }  )+$signed( { 2'b0,x191 } <<<3'd1 )+$signed( { 3'b0,x192 }<<<3'd2 )+$signed( { 2'b0,x193 } <<<3'd1 )+$signed( -{ 1'b0,x194 } )+$signed( { 1'b0,x195 }  )+$signed( { 3'b0,x196 }<<<3'd2 )+$signed( { 2'b0,x197 } <<<3'd1 )+$signed( -{ 2'b0,x198 }<<<3'd1 )+$signed( -{ 2'b0,x199 }<<<3'd1 )+$signed( -{ 3'b0,x200 }<<<3'd2)+$signed( -{ 3'b0,x201 }<<<3'd2)+$signed( -{ 2'b0,x202 }<<<3'd1 )+$signed( -{ 1'b0,x203 } )+$signed( { 2'b0,x204 } <<<3'd1 )+$signed( { 2'b0,x205 } <<<3'd1 )+$signed( -{ 1'b0,x206 } )+$signed( { 1'b0,x207 }  )+$signed( { 3'b0,x208 }<<<3'd2 )+$signed( { 1'b0,x210 }  )+$signed( -{ 1'b0,x211 } )+$signed( { 1'b0,x212 }  )+$signed( { 1'b0,x213 }  )+$signed( { 1'b0,x214 }  )+$signed( -{ 3'b0,x215 }<<<3'd2)+$signed( -{ 3'b0,x216 }<<<3'd2)+$signed( -{ 5'b0,x217 }<<<3'd4 )+$signed( { 3'b0,x218 }<<<3'd2 )+$signed( -{ 4'b0, x219 }<<<3'd3 )+$signed( -{ 2'b0,x220 }<<<3'd1 )+$signed( -{ 1'b0,x221 } )+$signed( { 3'b0,x222 }<<<3'd2 )+$signed( { 3'b0,x223 }<<<3'd2 )+$signed( { 1'b0,x224 }  )+$signed( { 2'b0,x225 } <<<3'd1 )+$signed( { 3'b0,x226 }<<<3'd2 )+$signed( -{ 2'b0,x228 }<<<3'd1 )+$signed( { 1'b0,x229 }  )+$signed( -{ 3'b0,x230 }<<<3'd2)+$signed( { 1'b0,x232 }  )+$signed( -{ 3'b0,x233 }<<<3'd2)+$signed( -{ 3'b0,x234 }<<<3'd2)+$signed( -{ 2'b0,x235 }<<<3'd1 )+$signed( -{ 4'b0, x237 }<<<3'd3 )+$signed( -{ 1'b0,x238 } )+$signed( { 1'b0,x239 }  )+$signed( { 3'b0,x240 }<<<3'd2 )+$signed( { 3'b0,x241 }<<<3'd2 )+$signed( { 1'b0,x242 }  )+$signed( { 1'b0,x243 }  )+$signed( { 2'b0,x244 } <<<3'd1 )+$signed( { 2'b0,x245 } <<<3'd1 )+$signed( -{ 2'b0,x246 }<<<3'd1 )+$signed( -{ 2'b0,x247 }<<<3'd1 )+$signed( { 2'b0,x248 } <<<3'd1 )+$signed( { 1'b0,x249 }  )+$signed( { 1'b0,x250 }  )+$signed( -{ 3'b0,x251 }<<<3'd2)+$signed( -{ 1'b0,x252 } )+$signed( { 2'b0,x254 } <<<3'd1 )+$signed( -{ 3'b0,x255 }<<<3'd2)+$signed( { 1'b0,x256 }  )+$signed( { 1'b0,x257 }  )+$signed( { 3'b0,x258 }<<<3'd2 )+$signed( -{ 1'b0,x259 } )+$signed( { 1'b0,x261 }  )+$signed( { 1'b0,x262 }  )+$signed( -{ 3'b0,x264 }<<<3'd2)+$signed( -{ 1'b0,x265 } )+$signed( -{ 1'b0,x266 } )+$signed( { 2'b0,x267 } <<<3'd1 )+$signed( { 2'b0,x268 } <<<3'd1 )+$signed( -{ 3'b0,x269 }<<<3'd2)+$signed( -{ 2'b0,x270 }<<<3'd1 )+$signed( -{ 1'b0,x271 } )+$signed( -{ 2'b0,x272 }<<<3'd1 )+$signed( -{ 3'b0,x273 }<<<3'd2)+$signed( -{ 3'b0,x274 }<<<3'd2)+$signed( -{ 1'b0,x275 } )+$signed( { 3'b0,x276 }<<<3'd2 )+$signed( { 3'b0,x277 }<<<3'd2 )+$signed( { 1'b0,x278 }  )+$signed( -{ 1'b0,x279 } )+$signed( { 3'b0,x280 }<<<3'd2 )+$signed( -{ 3'b0,x281 }<<<3'd2)+$signed( -{ 1'b0,x282 } )+$signed( -{ 2'b0,x283 }<<<3'd1 )+$signed( { 2'b0,x284 } <<<3'd1 )+$signed( { 1'b0,x285 }  )+$signed( -{ 2'b0,x286 }<<<3'd1 )+$signed( -{ 2'b0,x287 }<<<3'd1 )+$signed( -{ 3'b0,x288 }<<<3'd2)+$signed( { 2'b0,x289 } <<<3'd1 )+$signed( { 1'b0,x290 }  )+$signed( -{ 1'b0,x291 } )+$signed( -{ 3'b0,x292 }<<<3'd2)+$signed( -{ 2'b0,x293 }<<<3'd1 )+$signed( -{ 1'b0,x294 } )+$signed( { 2'b0,x295 } <<<3'd1 )+$signed( { 1'b0,x296 }  )+$signed( -{ 2'b0,x297 }<<<3'd1 )+$signed( -{ 2'b0,x298 }<<<3'd1 )+$signed( -{ 4'b0, x299 }<<<3'd3 )+$signed( { 2'b0,x300 } <<<3'd1 )+$signed( { 2'b0,x302 } <<<3'd1 )+$signed( -{ 2'b0,x303 }<<<3'd1 )+$signed( -{ 3'b0,x304 }<<<3'd2)+$signed( -{ 3'b0,x305 }<<<3'd2)+$signed( -{ 2'b0,x306 }<<<3'd1 )+$signed( -{ 1'b0,x307 } )+$signed( { 1'b0,x308 }  )+$signed( { 3'b0,x309 }<<<3'd2 )+$signed( { 2'b0,x310 } <<<3'd1 )+$signed( { 1'b0,x311 }  )+$signed( -{ 3'b0,x312 }<<<3'd2)+$signed( { 1'b0,x313 }  )+$signed( -{ 2'b0,x314 }<<<3'd1 )+$signed( -{ 1'b0,x315 } )+$signed( -{ 2'b0,x316 }<<<3'd1 )+$signed( -{ 1'b0,x317 } )+$signed( { 2'b0,x318 } <<<3'd1 )+$signed( -{ 1'b0,x319 } )+$signed( -{ 1'b0,x320 } )+$signed( { 2'b0,x321 } <<<3'd1 )+$signed( { 1'b0,x323 }  )+$signed( -{ 1'b0,x324 } )+$signed( -{ 3'b0,x325 }<<<3'd2)+$signed( { 1'b0,x326 }  )+$signed( -{ 1'b0,x327 } )+$signed( { 2'b0,x328 } <<<3'd1 )+$signed( { 1'b0,x329 }  )+$signed( -{ 1'b0,x330 } )+$signed( -{ 2'b0,x331 }<<<3'd1 )+$signed( -{ 3'b0,x332 }<<<3'd2)+$signed( -{ 2'b0,x333 }<<<3'd1 )+$signed( { 3'b0,x334 }<<<3'd2 )+$signed( { 2'b0,x336 } <<<3'd1 )+$signed( -{ 1'b0,x337 } )+$signed( -{ 2'b0,x338 }<<<3'd1 )+$signed( { 1'b0,x339 }  )+$signed( -{ 1'b0,x340 } )+$signed( { 2'b0,x341 } <<<3'd1 )+$signed( -{ 3'b0,x343 }<<<3'd2)+$signed( -{ 4'b0, x344 }<<<3'd3 )+$signed( -{ 2'b0,x345 }<<<3'd1 )+$signed( -{ 2'b0,x346 }<<<3'd1 )+$signed( { 3'b0,x347 }<<<3'd2 )+$signed( { 1'b0,x348 }  )+$signed( { 2'b0,x349 } <<<3'd1 )+$signed( { 1'b0,x350 }  )+$signed( -{ 5'b0,x351 }<<<3'd4 )+$signed( -{ 1'b0,x352 } )+$signed( { 2'b0,x353 } <<<3'd1 )+$signed( { 2'b0,x354 } <<<3'd1 )+$signed( -{ 1'b0,x355 } )+$signed( -{ 3'b0,x356 }<<<3'd2)+$signed( -{ 3'b0,x357 }<<<3'd2)+$signed( -{ 2'b0,x358 }<<<3'd1 )+$signed( -{ 1'b0,x359 } )+$signed( { 2'b0,x360 } <<<3'd1 )+$signed( { 1'b0,x361 }  )+$signed( { 2'b0,x362 } <<<3'd1 )+$signed( { 1'b0,x363 }  )+$signed( { 2'b0,x364 } <<<3'd1 )+$signed( -{ 2'b0,x365 }<<<3'd1 )+$signed( -{ 1'b0,x366 } )+$signed( -{ 2'b0,x368 }<<<3'd1 )+$signed( -{ 2'b0,x369 }<<<3'd1 )+$signed( { 1'b0,x370 }  )+$signed( -{ 3'b0,x371 }<<<3'd2)+$signed( { 1'b0,x372 }  )+$signed( { 2'b0,x373 } <<<3'd1 )+$signed( { 3'b0,x374 }<<<3'd2 )+$signed( -{ 2'b0,x375 }<<<3'd1 )+$signed( -{ 2'b0,x376 }<<<3'd1 )+$signed( -{ 2'b0,x377 }<<<3'd1 )+$signed( -{ 2'b0,x378 }<<<3'd1 )+$signed( -{ 3'b0,x379 }<<<3'd2)+$signed( { 2'b0,x380 } <<<3'd1 )+$signed( -{ 3'b0,x381 }<<<3'd2)+$signed( -{ 2'b0,x382 }<<<3'd1 )+$signed( -{ 2'b0,x383 }<<<3'd1 )+$signed( -{ 2'b0,x384 }<<<3'd1 )+$signed( { 2'b0,x385 } <<<3'd1 )+$signed( { 2'b0,x386 } <<<3'd1 )+$signed( { 3'b0,x387 }<<<3'd2 )+$signed( { 3'b0,x388 }<<<3'd2 )+$signed( { 1'b0,x389 }  )+$signed( { 2'b0,x391 } <<<3'd1 )+$signed( { 1'b0,x393 }  )+$signed( { 1'b0,x394 }  )+$signed( { 1'b0,x395 }  )+$signed( -{ 2'b0,x396 }<<<3'd1 )+$signed( { 1'b0,x397 }  )+$signed( { 2'b0,x398 } <<<3'd1 )+$signed( { 3'b0,x399 }<<<3'd2 )+$signed( { 1'b0,x400 }  )+$signed( -{ 2'b0,x402 }<<<3'd1 )+$signed( -{ 4'b0, x403 }<<<3'd3 )+$signed( -{ 2'b0,x404 }<<<3'd1 )+$signed( { 3'b0,x406 }<<<3'd2 )+$signed( -{ 2'b0,x407 }<<<3'd1 )+$signed( -{ 4'b0, x408 }<<<3'd3 )+$signed( -{ 1'b0,x409 } )+$signed( -{ 3'b0,x410 }<<<3'd2)+$signed( -{ 1'b0,x411 } )+$signed( { 3'b0,x412 }<<<3'd2 )+$signed( -{ 1'b0,x413 } )+$signed( { 3'b0,x414 }<<<3'd2 )+$signed( { 3'b0,x415 }<<<3'd2 )+$signed( -{ 3'b0,x417 }<<<3'd2)+$signed( -{ 3'b0,x418 }<<<3'd2)+$signed( { 1'b0,x419 }  )+$signed( { 2'b0,x420 } <<<3'd1 )+$signed( -{ 3'b0,x421 }<<<3'd2)+$signed( -{ 3'b0,x422 }<<<3'd2)+$signed( { 2'b0,x423 } <<<3'd1 )+$signed( { 3'b0,x424 }<<<3'd2 )+$signed( { 1'b0,x425 }  )+$signed( { 2'b0,x427 } <<<3'd1 )+$signed( { 1'b0,x428 }  )+$signed( -{ 4'b0, x429 }<<<3'd3 )+$signed( { 2'b0,x430 } <<<3'd1 )+$signed( { 3'b0,x432 }<<<3'd2 )+$signed( -{ 3'b0,x433 }<<<3'd2)+$signed( -{ 1'b0,x434 } )+$signed( -{ 3'b0,x435 }<<<3'd2)+$signed( -{ 3'b0,x436 }<<<3'd2)+$signed( { 3'b0,x439 }<<<3'd2 )+$signed( { 2'b0,x441 } <<<3'd1 )+$signed( -{ 3'b0,x442 }<<<3'd2)+$signed( { 2'b0,x443 } <<<3'd1 )+$signed( { 2'b0,x444 } <<<3'd1 )+$signed( { 2'b0,x445 } <<<3'd1 )+$signed( -{ 1'b0,x446 } )+$signed( -{ 3'b0,x447 }<<<3'd2)+$signed( -{ 3'b0,x448 }<<<3'd2)+$signed( -{ 1'b0,x449 } )+$signed( { 3'b0,x451 }<<<3'd2 )+$signed( -{ 2'b0,x452 }<<<3'd1 )+$signed( { 2'b0,x453 } <<<3'd1 )+$signed( -{ 1'b0,x454 } )+$signed( -{ 4'b0, x455 }<<<3'd3 )+$signed( -{ 3'b0,x456 }<<<3'd2)+$signed( { 1'b0,x457 }  )+$signed( { 3'b0,x458 }<<<3'd2 )+$signed( { 3'b0,x459 }<<<3'd2 )+$signed( -{ 3'b0,x461 }<<<3'd2)+$signed( -{ 2'b0,x462 }<<<3'd1 )+$signed( { 3'b0,x464 }<<<3'd2 )+$signed( { 3'b0,x465 }<<<3'd2 )+$signed( { 3'b0,x466 }<<<3'd2 )+$signed( { 2'b0,x467 } <<<3'd1 )+$signed( -{ 1'b0,x468 } )+$signed( -{ 2'b0,x469 }<<<3'd1 )+$signed( -{ 3'b0,x470 }<<<3'd2)+$signed( { 3'b0,x471 }<<<3'd2 )+$signed( -{ 2'b0,x472 }<<<3'd1 )+$signed( -{ 2'b0,x473 }<<<3'd1 )+$signed( -{ 2'b0,x474 }<<<3'd1 )+$signed( -{ 3'b0,x475 }<<<3'd2)+$signed( { 1'b0,x476 }  )+$signed( { 3'b0,x477 }<<<3'd2 )+$signed( { 2'b0,x478 } <<<3'd1 )+$signed( { 2'b0,x479 } <<<3'd1 )+$signed( -{ 3'b0,x481 }<<<3'd2)+$signed( -{ 1'b0,x482 } )+$signed( -{ 2'b0,x483 }<<<3'd1 )+$signed( { 3'b0,x484 }<<<3'd2 )+$signed( -{ 3'b0,x485 }<<<3'd2)+$signed( { 2'b0,x486 } <<<3'd1 )+$signed( -{ 3'b0,x487 }<<<3'd2)+$signed( -{ 1'b0,x488 } )+$signed( { 3'b0,x490 }<<<3'd2 )+$signed( { 1'b0,x491 }  )+$signed( { 1'b0,x492 }  )+$signed( { 1'b0,x493 }  )+$signed( -{ 3'b0,x494 }<<<3'd2)+$signed(13'd72);
assign y19=temp_y[19][13] ==1'b1 ? 6'd0 :  
    temp_y[19][10] ==1'b1 ? 6'd63 : 
    temp_y[19][3]==1'b1 ? temp_y[19][9:4]+1'b1 : temp_y[19][9:4];
endmodule