module Dense1(
input [4:0] x0 ,
input [4:0] x1 ,
input [4:0] x2 ,
input [4:0] x3 ,
input [4:0] x4 ,
input [4:0] x5 ,
input [4:0] x6 ,
input [4:0] x7 ,
input [4:0] x8 ,
input [4:0] x9 ,
input [4:0] x10 ,
input [4:0] x11 ,
input [4:0] x12 ,
input [4:0] x13 ,
input [4:0] x14 ,
input [4:0] x15 ,
input [4:0] x16 ,
input [4:0] x17 ,
input [4:0] x18 ,
input [4:0] x19 ,
input [4:0] x20 ,
input [4:0] x21 ,
input [4:0] x22 ,
input [4:0] x23 ,
input [4:0] x24 ,
input [4:0] x25 ,
input [4:0] x26 ,
input [4:0] x27 ,
input [4:0] x28 ,
input [4:0] x29 ,
input [4:0] x30 ,
input [4:0] x31 ,
input [4:0] x32 ,
input [4:0] x33 ,
input [4:0] x34 ,
input [4:0] x35 ,
input [4:0] x36 ,
input [4:0] x37 ,
input [4:0] x38 ,
input [4:0] x39 ,
input [4:0] x40 ,
input [4:0] x41 ,
input [4:0] x42 ,
input [4:0] x43 ,
input [4:0] x44 ,
input [4:0] x45 ,
input [4:0] x46 ,
input [4:0] x47 ,
input [4:0] x48 ,
input [4:0] x49 ,
input [4:0] x50 ,
input [4:0] x51 ,
input [4:0] x52 ,
input [4:0] x53 ,
input [4:0] x54 ,
input [4:0] x55 ,
input [4:0] x56 ,
input [4:0] x57 ,
input [4:0] x58 ,
input [4:0] x59 ,
input [4:0] x60 ,
input [4:0] x61 ,
input [4:0] x62 ,
input [4:0] x63 ,
input [4:0] x64 ,
input [4:0] x65 ,
input [4:0] x66 ,
input [4:0] x67 ,
input [4:0] x68 ,
input [4:0] x69 ,
input [4:0] x70 ,
input [4:0] x71 ,
input [4:0] x72 ,
input [4:0] x73 ,
input [4:0] x74 ,
input [4:0] x75 ,
input [4:0] x76 ,
input [4:0] x77 ,
input [4:0] x78 ,
input [4:0] x79 ,
input [4:0] x80 ,
input [4:0] x81 ,
input [4:0] x82 ,
input [4:0] x83 ,
input [4:0] x84 ,
input [4:0] x85 ,
input [4:0] x86 ,
input [4:0] x87 ,
input [4:0] x88 ,
input [4:0] x89 ,
input [4:0] x90 ,
input [4:0] x91 ,
input [4:0] x92 ,
input [4:0] x93 ,
input [4:0] x94 ,
input [4:0] x95 ,
input [4:0] x96 ,
input [4:0] x97 ,
input [4:0] x98 ,
input [4:0] x99 ,
input [4:0] x100 ,
input [4:0] x101 ,
input [4:0] x102 ,
input [4:0] x103 ,
input [4:0] x104 ,
input [4:0] x105 ,
input [4:0] x106 ,
input [4:0] x107 ,
input [4:0] x108 ,
input [4:0] x109 ,
input [4:0] x110 ,
input [4:0] x111 ,
input [4:0] x112 ,
input [4:0] x113 ,
input [4:0] x114 ,
input [4:0] x115 ,
input [4:0] x116 ,
input [4:0] x117 ,
input [4:0] x118 ,
input [4:0] x119 ,
input [4:0] x120 ,
input [4:0] x121 ,
input [4:0] x122 ,
input [4:0] x123 ,
input [4:0] x124 ,
input [4:0] x125 ,
input [4:0] x126 ,
input [4:0] x127 ,
input [4:0] x128 ,
input [4:0] x129 ,
input [4:0] x130 ,
input [4:0] x131 ,
input [4:0] x132 ,
input [4:0] x133 ,
input [4:0] x134 ,
input [4:0] x135 ,
input [4:0] x136 ,
input [4:0] x137 ,
input [4:0] x138 ,
input [4:0] x139 ,
input [4:0] x140 ,
input [4:0] x141 ,
input [4:0] x142 ,
input [4:0] x143 ,
input [4:0] x144 ,
input [4:0] x145 ,
input [4:0] x146 ,
input [4:0] x147 ,
input [4:0] x148 ,
input [4:0] x149 ,
input [4:0] x150 ,
input [4:0] x151 ,
input [4:0] x152 ,
input [4:0] x153 ,
input [4:0] x154 ,
input [4:0] x155 ,
input [4:0] x156 ,
input [4:0] x157 ,
input [4:0] x158 ,
input [4:0] x159 ,
input [4:0] x160 ,
input [4:0] x161 ,
input [4:0] x162 ,
input [4:0] x163 ,
input [4:0] x164 ,
input [4:0] x165 ,
input [4:0] x166 ,
input [4:0] x167 ,
input [4:0] x168 ,
input [4:0] x169 ,
input [4:0] x170 ,
input [4:0] x171 ,
input [4:0] x172 ,
input [4:0] x173 ,
input [4:0] x174 ,
input [4:0] x175 ,
input [4:0] x176 ,
input [4:0] x177 ,
input [4:0] x178 ,
input [4:0] x179 ,
input [4:0] x180 ,
input [4:0] x181 ,
input [4:0] x182 ,
input [4:0] x183 ,
input [4:0] x184 ,
input [4:0] x185 ,
input [4:0] x186 ,
input [4:0] x187 ,
input [4:0] x188 ,
input [4:0] x189 ,
input [4:0] x190 ,
input [4:0] x191 ,
input [4:0] x192 ,
input [4:0] x193 ,
input [4:0] x194 ,
input [4:0] x195 ,
input [4:0] x196 ,
input [4:0] x197 ,
input [4:0] x198 ,
input [4:0] x199 ,
input [4:0] x200 ,
input [4:0] x201 ,
input [4:0] x202 ,
input [4:0] x203 ,
input [4:0] x204 ,
input [4:0] x205 ,
input [4:0] x206 ,
input [4:0] x207 ,
input [4:0] x208 ,
input [4:0] x209 ,
input [4:0] x210 ,
input [4:0] x211 ,
input [4:0] x212 ,
input [4:0] x213 ,
input [4:0] x214 ,
input [4:0] x215 ,
input [4:0] x216 ,
input [4:0] x217 ,
input [4:0] x218 ,
input [4:0] x219 ,
input [4:0] x220 ,
input [4:0] x221 ,
input [4:0] x222 ,
input [4:0] x223 ,
input [4:0] x224 ,
input [4:0] x225 ,
input [4:0] x226 ,
input [4:0] x227 ,
input [4:0] x228 ,
input [4:0] x229 ,
input [4:0] x230 ,
input [4:0] x231 ,
input [4:0] x232 ,
input [4:0] x233 ,
input [4:0] x234 ,
input [4:0] x235 ,
input [4:0] x236 ,
input [4:0] x237 ,
input [4:0] x238 ,
input [4:0] x239 ,
input [4:0] x240 ,
input [4:0] x241 ,
input [4:0] x242 ,
input [4:0] x243 ,
input [4:0] x244 ,
input [4:0] x245 ,
input [4:0] x246 ,
input [4:0] x247 ,
input [4:0] x248 ,
input [4:0] x249 ,
input [4:0] x250 ,
input [4:0] x251 ,
input [4:0] x252 ,
input [4:0] x253 ,
input [4:0] x254 ,
input [4:0] x255 ,
input [4:0] x256 ,
input [4:0] x257 ,
input [4:0] x258 ,
input [4:0] x259 ,
input [4:0] x260 ,
input [4:0] x261 ,
input [4:0] x262 ,
input [4:0] x263 ,
input [4:0] x264 ,
input [4:0] x265 ,
input [4:0] x266 ,
input [4:0] x267 ,
input [4:0] x268 ,
input [4:0] x269 ,
input [4:0] x270 ,
input [4:0] x271 ,
input [4:0] x272 ,
input [4:0] x273 ,
input [4:0] x274 ,
input [4:0] x275 ,
input [4:0] x276 ,
input [4:0] x277 ,
input [4:0] x278 ,
input [4:0] x279 ,
input [4:0] x280 ,
input [4:0] x281 ,
input [4:0] x282 ,
input [4:0] x283 ,
input [4:0] x284 ,
input [4:0] x285 ,
input [4:0] x286 ,
input [4:0] x287 ,
input [4:0] x288 ,
input [4:0] x289 ,
input [4:0] x290 ,
input [4:0] x291 ,
input [4:0] x292 ,
input [4:0] x293 ,
input [4:0] x294 ,
input [4:0] x295 ,
input [4:0] x296 ,
input [4:0] x297 ,
input [4:0] x298 ,
input [4:0] x299 ,
input [4:0] x300 ,
input [4:0] x301 ,
input [4:0] x302 ,
input [4:0] x303 ,
input [4:0] x304 ,
input [4:0] x305 ,
input [4:0] x306 ,
input [4:0] x307 ,
input [4:0] x308 ,
input [4:0] x309 ,
input [4:0] x310 ,
input [4:0] x311 ,
input [4:0] x312 ,
input [4:0] x313 ,
input [4:0] x314 ,
input [4:0] x315 ,
input [4:0] x316 ,
input [4:0] x317 ,
input [4:0] x318 ,
input [4:0] x319 ,
input [4:0] x320 ,
input [4:0] x321 ,
input [4:0] x322 ,
input [4:0] x323 ,
input [4:0] x324 ,
input [4:0] x325 ,
input [4:0] x326 ,
input [4:0] x327 ,
input [4:0] x328 ,
input [4:0] x329 ,
input [4:0] x330 ,
input [4:0] x331 ,
input [4:0] x332 ,
input [4:0] x333 ,
input [4:0] x334 ,
input [4:0] x335 ,
input [4:0] x336 ,
input [4:0] x337 ,
input [4:0] x338 ,
input [4:0] x339 ,
input [4:0] x340 ,
input [4:0] x341 ,
input [4:0] x342 ,
input [4:0] x343 ,
input [4:0] x344 ,
input [4:0] x345 ,
input [4:0] x346 ,
input [4:0] x347 ,
input [4:0] x348 ,
input [4:0] x349 ,
input [4:0] x350 ,
input [4:0] x351 ,
input [4:0] x352 ,
input [4:0] x353 ,
input [4:0] x354 ,
input [4:0] x355 ,
input [4:0] x356 ,
input [4:0] x357 ,
input [4:0] x358 ,
input [4:0] x359 ,
input [4:0] x360 ,
input [4:0] x361 ,
input [4:0] x362 ,
input [4:0] x363 ,
input [4:0] x364 ,
input [4:0] x365 ,
input [4:0] x366 ,
input [4:0] x367 ,
input [4:0] x368 ,
input [4:0] x369 ,
input [4:0] x370 ,
input [4:0] x371 ,
input [4:0] x372 ,
input [4:0] x373 ,
input [4:0] x374 ,
input [4:0] x375 ,
input [4:0] x376 ,
input [4:0] x377 ,
input [4:0] x378 ,
input [4:0] x379 ,
input [4:0] x380 ,
input [4:0] x381 ,
input [4:0] x382 ,
input [4:0] x383 ,
input [4:0] x384 ,
input [4:0] x385 ,
input [4:0] x386 ,
input [4:0] x387 ,
input [4:0] x388 ,
input [4:0] x389 ,
input [4:0] x390 ,
input [4:0] x391 ,
input [4:0] x392 ,
input [4:0] x393 ,
input [4:0] x394 ,
input [4:0] x395 ,
input [4:0] x396 ,
input [4:0] x397 ,
input [4:0] x398 ,
input [4:0] x399 ,
input [4:0] x400 ,
input [4:0] x401 ,
input [4:0] x402 ,
input [4:0] x403 ,
input [4:0] x404 ,
input [4:0] x405 ,
input [4:0] x406 ,
input [4:0] x407 ,
input [4:0] x408 ,
input [4:0] x409 ,
input [4:0] x410 ,
input [4:0] x411 ,
input [4:0] x412 ,
input [4:0] x413 ,
input [4:0] x414 ,
input [4:0] x415 ,
input [4:0] x416 ,
input [4:0] x417 ,
input [4:0] x418 ,
input [4:0] x419 ,
input [4:0] x420 ,
input [4:0] x421 ,
input [4:0] x422 ,
input [4:0] x423 ,
input [4:0] x424 ,
input [4:0] x425 ,
input [4:0] x426 ,
input [4:0] x427 ,
input [4:0] x428 ,
input [4:0] x429 ,
input [4:0] x430 ,
input [4:0] x431 ,
input [4:0] x432 ,
input [4:0] x433 ,
input [4:0] x434 ,
input [4:0] x435 ,
input [4:0] x436 ,
input [4:0] x437 ,
input [4:0] x438 ,
input [4:0] x439 ,
input [4:0] x440 ,
input [4:0] x441 ,
input [4:0] x442 ,
input [4:0] x443 ,
input [4:0] x444 ,
input [4:0] x445 ,
input [4:0] x446 ,
input [4:0] x447 ,
input [4:0] x448 ,
input [4:0] x449 ,
input [4:0] x450 ,
input [4:0] x451 ,
input [4:0] x452 ,
input [4:0] x453 ,
input [4:0] x454 ,
input [4:0] x455 ,
input [4:0] x456 ,
input [4:0] x457 ,
input [4:0] x458 ,
input [4:0] x459 ,
input [4:0] x460 ,
input [4:0] x461 ,
input [4:0] x462 ,
input [4:0] x463 ,
input [4:0] x464 ,
input [4:0] x465 ,
input [4:0] x466 ,
input [4:0] x467 ,
input [4:0] x468 ,
input [4:0] x469 ,
input [4:0] x470 ,
input [4:0] x471 ,
input [4:0] x472 ,
input [4:0] x473 ,
input [4:0] x474 ,
input [4:0] x475 ,
input [4:0] x476 ,
input [4:0] x477 ,
input [4:0] x478 ,
input [4:0] x479 ,
input [4:0] x480 ,
input [4:0] x481 ,
input [4:0] x482 ,
input [4:0] x483 ,
input [4:0] x484 ,
input [4:0] x485 ,
input [4:0] x486 ,
input [4:0] x487 ,
input [4:0] x488 ,
input [4:0] x489 ,
input [4:0] x490 ,
input [4:0] x491 ,
input [4:0] x492 ,
input [4:0] x493 ,
input [4:0] x494 ,
input [4:0] x495 ,
output [5:0] y0 ,
output [5:0] y1 ,
output [5:0] y2 ,
output [5:0] y3 ,
output [5:0] y4 ,
output [5:0] y5 ,
output [5:0] y6 ,
output [5:0] y7 ,
output [5:0] y8 ,
output [5:0] y9 ,
output [5:0] y10 ,
output [5:0] y11 ,
output [5:0] y12 ,
output [5:0] y13 ,
output [5:0] y14 ,
output [5:0] y15 ,
output [5:0] y16 ,
output [5:0] y17 ,
output [5:0] y18 ,
output [5:0] y19 
);
wire [13:0] sharing0;
wire [13:0] sharing1;
wire [13:0] sharing2;
wire [13:0] sharing3;
wire [13:0] sharing4;
wire [13:0] sharing5;
wire [13:0] sharing6;
wire [13:0] sharing7;
wire [13:0] sharing8;
wire [13:0] sharing9;
wire [13:0] sharing10;
wire [13:0] sharing11;
wire [13:0] sharing12;
wire [13:0] sharing13;
wire [13:0] sharing14;
wire [13:0] sharing15;
wire [13:0] sharing16;
wire [13:0] sharing17;
wire [13:0] sharing18;
wire [13:0] sharing19;
wire [13:0] sharing20;
wire [13:0] sharing21;
wire [13:0] sharing22;
wire [13:0] sharing23;
wire [13:0] sharing24;
wire [13:0] sharing25;
wire [13:0] sharing26;
wire [13:0] sharing27;
wire [13:0] sharing28;
wire [13:0] sharing29;
wire [13:0] sharing30;
wire [13:0] sharing31;
wire [13:0] sharing32;
wire [13:0] sharing33;
wire [13:0] sharing34;
wire [13:0] sharing35;
wire [13:0] sharing36;
wire [13:0] sharing37;
wire [13:0] sharing38;
wire [13:0] sharing39;
wire [13:0] sharing40;
wire [13:0] sharing41;
wire [13:0] sharing42;
wire [13:0] sharing43;
wire [13:0] sharing44;
wire [13:0] sharing45;
wire [13:0] sharing46;
wire [13:0] sharing47;
wire [13:0] sharing48;
wire [13:0] sharing49;
wire [13:0] sharing50;
wire [13:0] sharing51;
wire [13:0] sharing52;
wire [13:0] sharing53;
wire [13:0] sharing54;
wire [13:0] sharing55;
wire [13:0] sharing56;
wire [13:0] sharing57;
wire [13:0] sharing58;
wire [13:0] sharing59;
wire [13:0] sharing60;
wire [13:0] sharing61;
wire [13:0] sharing62;
wire [13:0] sharing63;
wire [13:0] sharing64;
wire [13:0] sharing65;
wire [13:0] sharing66;
wire [13:0] sharing67;
wire [13:0] sharing68;
wire [13:0] sharing69;
wire [13:0] sharing70;
wire [13:0] sharing71;
wire [13:0] sharing72;
wire [13:0] sharing73;
wire [13:0] sharing74;
wire [13:0] sharing75;
wire [13:0] sharing76;
wire [13:0] sharing77;
wire [13:0] sharing78;
wire [13:0] sharing79;
wire [13:0] sharing80;
wire [13:0] sharing81;
wire [13:0] sharing82;
wire [13:0] sharing83;
wire [13:0] sharing84;
wire [13:0] sharing85;
wire [13:0] sharing86;
wire [13:0] sharing87;
wire [13:0] sharing88;
wire [13:0] sharing89;
wire [13:0] sharing90;
wire [13:0] sharing91;
wire [13:0] sharing92;
wire [13:0] sharing93;
wire [13:0] sharing94;
wire [13:0] sharing95;
wire [13:0] sharing96;
wire [13:0] sharing97;
wire [13:0] sharing98;
wire [13:0] sharing99;
wire [13:0] sharing100;
wire [13:0] sharing101;
wire [13:0] sharing102;
wire [13:0] sharing103;
wire [13:0] sharing104;
wire [13:0] sharing105;
wire [13:0] sharing106;
wire [13:0] sharing107;
wire [13:0] sharing108;
wire [13:0] sharing109;
wire [13:0] sharing110;
wire [13:0] sharing111;
wire [13:0] sharing112;
wire [13:0] sharing113;
wire [13:0] sharing114;
wire [13:0] sharing115;
wire [13:0] sharing116;
wire [13:0] sharing117;
wire [13:0] sharing118;
wire [13:0] sharing119;
wire [13:0] sharing120;
wire [13:0] sharing121;
wire [13:0] sharing122;
wire [13:0] sharing123;
wire [13:0] sharing124;
wire [13:0] sharing125;
wire [13:0] sharing126;
wire [13:0] sharing127;
wire [13:0] sharing128;
wire [13:0] sharing129;
wire [13:0] sharing130;
wire [13:0] sharing131;
wire [13:0] sharing132;
wire [13:0] sharing133;
wire [13:0] sharing134;
wire [13:0] sharing135;
wire [13:0] sharing136;
wire [13:0] sharing137;
wire [13:0] sharing138;
wire [13:0] sharing139;
wire [13:0] sharing140;
wire [13:0] sharing141;
wire [13:0] sharing142;
wire [13:0] sharing143;
wire [13:0] sharing144;
wire [13:0] sharing145;
wire [13:0] sharing146;
wire [13:0] sharing147;
wire [13:0] sharing148;
wire [13:0] sharing149;
wire [13:0] sharing150;
wire [13:0] sharing151;
wire [13:0] sharing152;
wire [13:0] sharing153;
wire [13:0] sharing154;
wire [13:0] sharing155;
wire [13:0] sharing156;
wire [13:0] sharing157;
wire [13:0] sharing158;
wire [13:0] sharing159;
wire [13:0] sharing160;
wire [13:0] sharing161;
wire [13:0] sharing162;
wire [13:0] sharing163;
wire [13:0] sharing164;
wire [13:0] sharing165;
wire [13:0] sharing166;
wire [13:0] sharing167;
wire [13:0] sharing168;
wire [13:0] sharing169;
wire [13:0] sharing170;
wire [13:0] sharing171;
wire [13:0] sharing172;
wire [13:0] sharing173;
wire [13:0] sharing174;
wire [13:0] sharing175;
wire [13:0] sharing176;
wire [13:0] sharing177;
wire [13:0] sharing178;
wire [13:0] sharing179;
wire [13:0] sharing180;
wire [13:0] sharing181;
wire [13:0] sharing182;
wire [13:0] sharing183;
wire [13:0] sharing184;
wire [13:0] sharing185;
wire [13:0] sharing186;
wire [13:0] sharing187;
wire [13:0] sharing188;
wire [13:0] sharing189;
wire [13:0] sharing190;
wire [13:0] sharing191;
wire [13:0] sharing192;
wire [13:0] sharing193;
wire [13:0] sharing194;
wire [13:0] sharing195;
wire [13:0] sharing196;
wire [13:0] sharing197;
wire [13:0] sharing198;
wire [13:0] sharing199;
wire [13:0] sharing200;
wire [13:0] sharing201;
wire [13:0] sharing202;
wire [13:0] sharing203;
wire [13:0] sharing204;
wire [13:0] sharing205;
wire [13:0] sharing206;
wire [13:0] sharing207;
wire [13:0] sharing208;
wire [13:0] sharing209;
wire [13:0] sharing210;
wire [13:0] sharing211;
wire [13:0] sharing212;
wire [13:0] sharing213;
wire [13:0] sharing214;
wire [13:0] sharing215;
wire [13:0] sharing216;
wire [13:0] sharing217;
wire [13:0] sharing218;
wire [13:0] sharing219;
wire [13:0] sharing220;
wire [13:0] sharing221;
wire [13:0] sharing222;
wire [13:0] sharing223;
wire [13:0] sharing224;
wire [13:0] sharing225;
wire [13:0] sharing226;
wire [13:0] sharing227;
wire [13:0] sharing228;
wire [13:0] sharing229;
wire [13:0] sharing230;
wire [13:0] sharing231;
wire [13:0] sharing232;
wire [13:0] sharing233;
wire [13:0] sharing234;
wire [13:0] sharing235;
wire [13:0] sharing236;
wire [13:0] sharing237;
wire [13:0] sharing238;
wire [13:0] sharing239;
wire [13:0] sharing240;
wire [13:0] sharing241;
wire [13:0] sharing242;
wire [13:0] sharing243;
wire [13:0] sharing244;
wire [13:0] sharing245;
wire [13:0] sharing246;
wire [13:0] sharing247;
wire [13:0] sharing248;
wire [13:0] sharing249;
wire [13:0] sharing250;
wire [13:0] sharing251;
wire [13:0] sharing252;
wire [13:0] sharing253;
wire [13:0] sharing254;
wire [13:0] sharing255;
wire [13:0] sharing256;
wire [13:0] sharing257;
wire [13:0] sharing258;
wire [13:0] sharing259;
assign sharing0 = $signed(-{3'b0,x256}<<<3'd2)+$signed({2'b0,x416}<<<3'd1)+$signed({2'b0,x289}<<<3'd1)+$signed(-{3'b0,x226}<<<3'd2)+$signed({2'b0,x258}<<<3'd1)+$signed({3'b0,x355}<<<3'd2)+$signed(-{2'b0,x227}<<<3'd1)+$signed({1'b0,x35})+$signed(-{1'b0,x356})+$signed({3'b0,x421}<<<3'd2)+$signed(-{4'b0,x294}<<<3'd3)+$signed(-{3'b0,x454}<<<3'd2)+$signed({1'b0,x166})+$signed({2'b0,x231}<<<3'd1)+$signed({1'b0,x103})+$signed({3'b0,x392}<<<3'd2)+$signed({2'b0,x265}<<<3'd1)+$signed({2'b0,x457}<<<3'd1)+$signed({1'b0,x489})+$signed(-{1'b0,x233})+$signed(-{3'b0,x202}<<<3'd2)+$signed(-{2'b0,x234}<<<3'd1)+$signed(-{2'b0,x330}<<<3'd1)+$signed(-{1'b0,x427})+$signed({3'b0,x364}<<<3'd2)+$signed({2'b0,x268}<<<3'd1)+$signed(-{2'b0,x236}<<<3'd1)+$signed(-{2'b0,x428}<<<3'd1)+$signed({2'b0,x141}<<<3'd1)+$signed(-{2'b0,x333}<<<3'd1)+$signed({3'b0,x366}<<<3'd2)+$signed({2'b0,x110}<<<3'd1)+$signed(-{3'b0,x238}<<<3'd2)+$signed(-{3'b0,x271}<<<3'd2)+$signed({1'b0,x336})+$signed(-{4'b0,x337}<<<3'd3)+$signed({2'b0,x178}<<<3'd1)+$signed({1'b0,x210})+$signed(-{4'b0,x467}<<<3'd3)+$signed({3'b0,x115}<<<3'd2)+$signed(-{3'b0,x372}<<<3'd2)+$signed({2'b0,x276}<<<3'd1)+$signed(-{2'b0,x116}<<<3'd1)+$signed({3'b0,x21}<<<3'd2)+$signed(-{1'b0,x405})+$signed({3'b0,x118}<<<3'd2)+$signed({3'b0,x470}<<<3'd2)+$signed({3'b0,x471}<<<3'd2)+$signed({2'b0,x87}<<<3'd1)+$signed({1'b0,x247})+$signed(-{3'b0,x216}<<<3'd2)+$signed(-{3'b0,x376}<<<3'd2)+$signed(-{1'b0,x185})+$signed({2'b0,x90}<<<3'd1)+$signed({1'b0,x314})+$signed({3'b0,x347}<<<3'd2)+$signed({2'b0,x475}<<<3'd1)+$signed(-{2'b0,x59}<<<3'd1)+$signed(-{2'b0,x123}<<<3'd1)+$signed(-{3'b0,x92}<<<3'd2)+$signed(-{3'b0,x476}<<<3'd2)+$signed({1'b0,x412})+$signed(-{4'b0,x253}<<<3'd3)+$signed({3'b0,x93}<<<3'd2)+$signed(-{2'b0,x317}<<<3'd1)+$signed(-{3'b0,x286}<<<3'd2)+$signed({1'b0,x414})+$signed({2'b0,x159}<<<3'd1);
assign sharing1 = $signed({1'b0,x95})+$signed(-{1'b0,x162})+$signed({3'b0,x163}<<<3'd2)+$signed({2'b0,x419}<<<3'd1)+$signed(-{2'b0,x195}<<<3'd1)+$signed({3'b0,x260}<<<3'd2)+$signed({3'b0,x357}<<<3'd2)+$signed({3'b0,x133}<<<3'd2)+$signed({2'b0,x39}<<<3'd1)+$signed(-{3'b0,x40}<<<3'd2)+$signed({2'b0,x360}<<<3'd1)+$signed({1'b0,x72})+$signed(-{3'b0,x415}<<<3'd2)+$signed({1'b0,x425})+$signed(-{3'b0,x458}<<<3'd2)+$signed(-{3'b0,x426}<<<3'd2)+$signed({2'b0,x171}<<<3'd1)+$signed({2'b0,x203}<<<3'd1)+$signed({2'b0,x301}<<<3'd1)+$signed({3'b0,x207}<<<3'd2)+$signed({3'b0,x144}<<<3'd2)+$signed(-{3'b0,x112}<<<3'd2)+$signed(-{3'b0,x369}<<<3'd2)+$signed(-{2'b0,x401}<<<3'd1)+$signed({2'b0,x114}<<<3'd1)+$signed(-{2'b0,x466}<<<3'd1)+$signed(-{1'b0,x82})+$signed({3'b0,x243}<<<3'd2)+$signed({3'b0,x371}<<<3'd2)+$signed(-{1'b0,x434})+$signed(-{3'b0,x84}<<<3'd2)+$signed(-{3'b0,x148}<<<3'd2)+$signed(-{2'b0,x404}<<<3'd1)+$signed({2'b0,x469}<<<3'd1)+$signed({2'b0,x54}<<<3'd1)+$signed(-{2'b0,x310}<<<3'd1)+$signed({2'b0,x375}<<<3'd1)+$signed({3'b0,x88}<<<3'd2)+$signed({3'b0,x312}<<<3'd2)+$signed({1'b0,x153})+$signed({2'b0,x346}<<<3'd1)+$signed(-{2'b0,x58}<<<3'd1)+$signed({3'b0,x219}<<<3'd2)+$signed(-{3'b0,x27}<<<3'd2)+$signed(-{3'b0,x251}<<<3'd2)+$signed({3'b0,x316}<<<3'd2)+$signed({2'b0,x444}<<<3'd1)+$signed(-{3'b0,x252}<<<3'd2)+$signed(-{2'b0,x28}<<<3'd1)+$signed(-{3'b0,x445}<<<3'd2)+$signed({2'b0,x125}<<<3'd1)+$signed({2'b0,x157}<<<3'd1)+$signed(-{1'b0,x446})+$signed({3'b0,x479}<<<3'd2)+$signed({1'b0,x31});
assign sharing2 = $signed(-{3'b0,x448}<<<3'd2)+$signed(-{1'b0,x128})+$signed(-{3'b0,x193}<<<3'd2)+$signed({3'b0,x450}<<<3'd2)+$signed({3'b0,x483}<<<3'd2)+$signed(-{3'b0,x196}<<<3'd2)+$signed({2'b0,x36}<<<3'd1)+$signed(-{2'b0,x228}<<<3'd1)+$signed(-{1'b0,x4})+$signed(-{2'b0,x260}<<<3'd1)+$signed(-{3'b0,x133}<<<3'd2)+$signed(-{1'b0,x261})+$signed(-{1'b0,x5})+$signed({3'b0,x454}<<<3'd2)+$signed(-{2'b0,x70}<<<3'd1)+$signed(-{1'b0,x255})+$signed({2'b0,x7}<<<3'd1)+$signed({1'b0,x263})+$signed(-{2'b0,x199}<<<3'd1)+$signed(-{1'b0,x359})+$signed({3'b0,x201}<<<3'd2)+$signed(-{3'b0,x202}<<<3'd2)+$signed(-{2'b0,x426}<<<3'd1)+$signed({3'b0,x107}<<<3'd2)+$signed(-{3'b0,x299}<<<3'd2)+$signed(-{3'b0,x363}<<<3'd2)+$signed({3'b0,x429}<<<3'd2)+$signed(-{1'b0,x173})+$signed(-{3'b0,x366}<<<3'd2)+$signed(-{3'b0,x302}<<<3'd2)+$signed({1'b0,x110})+$signed(-{4'b0,x143}<<<3'd3)+$signed({3'b0,x431}<<<3'd2)+$signed(-{1'b0,x47})+$signed(-{2'b0,x368}<<<3'd1)+$signed(-{2'b0,x464}<<<3'd1)+$signed(-{2'b0,x179}<<<3'd1)+$signed(-{1'b0,x19})+$signed({3'b0,x340}<<<3'd2)+$signed({3'b0,x468}<<<3'd2)+$signed(-{3'b0,x116}<<<3'd2)+$signed({2'b0,x245}<<<3'd1)+$signed({3'b0,x214}<<<3'd2)+$signed({2'b0,x470}<<<3'd1)+$signed(-{2'b0,x406}<<<3'd1)+$signed(-{1'b0,x22})+$signed({3'b0,x183}<<<3'd2)+$signed(-{2'b0,x23}<<<3'd1)+$signed({3'b0,x184}<<<3'd2)+$signed({2'b0,x56}<<<3'd1)+$signed(-{2'b0,x376}<<<3'd1)+$signed({3'b0,x378}<<<3'd2)+$signed(-{3'b0,x154}<<<3'd2)+$signed(-{3'b0,x250}<<<3'd2)+$signed(-{3'b0,x444}<<<3'd2)+$signed({2'b0,x60}<<<3'd1)+$signed(-{2'b0,x348}<<<3'd1)+$signed(-{1'b0,x286})+$signed({3'b0,x159}<<<3'd2)+$signed(-{1'b0,x31});
assign sharing3 = $signed({3'b0,x416}<<<3'd2)+$signed({3'b0,x225}<<<3'd2)+$signed(-{3'b0,x98}<<<3'd2)+$signed(-{3'b0,x322}<<<3'd2)+$signed({3'b0,x163}<<<3'd2)+$signed(-{3'b0,x419}<<<3'd2)+$signed(-{2'b0,x227}<<<3'd1)+$signed(-{3'b0,x3}<<<3'd2)+$signed({1'b0,x101})+$signed({1'b0,x326})+$signed({3'b0,x392}<<<3'd2)+$signed(-{2'b0,x424}<<<3'd1)+$signed({1'b0,x40})+$signed(-{3'b0,x393}<<<3'd2)+$signed({3'b0,x234}<<<3'd2)+$signed({3'b0,x298}<<<3'd2)+$signed({3'b0,x330}<<<3'd2)+$signed(-{3'b0,x394}<<<3'd2)+$signed({3'b0,x171}<<<3'd2)+$signed(-{3'b0,x491}<<<3'd2)+$signed({3'b0,x236}<<<3'd2)+$signed(-{1'b0,x108})+$signed({4'b0,x461}<<<3'd3)+$signed({3'b0,x365}<<<3'd2)+$signed({3'b0,x430}<<<3'd2)+$signed({3'b0,x238}<<<3'd2)+$signed(-{3'b0,x462}<<<3'd2)+$signed({2'b0,x48}<<<3'd1)+$signed({1'b0,x336})+$signed({3'b0,x401}<<<3'd2)+$signed(-{2'b0,x242}<<<3'd1)+$signed(-{1'b0,x306})+$signed({3'b0,x339}<<<3'd2)+$signed({2'b0,x243}<<<3'd1)+$signed({3'b0,x371}<<<3'd2)+$signed({3'b0,x403}<<<3'd2)+$signed(-{3'b0,x467}<<<3'd2)+$signed({2'b0,x148}<<<3'd1)+$signed(-{3'b0,x341}<<<3'd2)+$signed({3'b0,x150}<<<3'd2)+$signed({3'b0,x438}<<<3'd2)+$signed({3'b0,x439}<<<3'd2)+$signed(-{3'b0,x215}<<<3'd2)+$signed({1'b0,x407})+$signed({4'b0,x120}<<<3'd3)+$signed({3'b0,x472}<<<3'd2)+$signed(-{2'b0,x151}<<<3'd1)+$signed(-{2'b0,x88}<<<3'd1)+$signed({3'b0,x121}<<<3'd2)+$signed({2'b0,x441}<<<3'd1)+$signed(-{3'b0,x186}<<<3'd2)+$signed({1'b0,x314})+$signed({3'b0,x411}<<<3'd2)+$signed({2'b0,x91}<<<3'd1)+$signed(-{3'b0,x251}<<<3'd2)+$signed(-{2'b0,x379}<<<3'd1)+$signed({1'b0,x124})+$signed({1'b0,x252})+$signed(-{1'b0,x380})+$signed(-{2'b0,x445}<<<3'd1)+$signed(-{3'b0,x222}<<<3'd2)+$signed({2'b0,x62}<<<3'd1)+$signed(-{1'b0,x126})+$signed(-{3'b0,x287}<<<3'd2)+$signed(-{1'b0,x447});
assign sharing4 = $signed({3'b0,x96}<<<3'd2)+$signed({2'b0,x352}<<<3'd1)+$signed({1'b0,x480})+$signed({3'b0,x385}<<<3'd2)+$signed(-{2'b0,x193}<<<3'd1)+$signed({1'b0,x289})+$signed(-{3'b0,x386}<<<3'd2)+$signed({3'b0,x387}<<<3'd2)+$signed(-{1'b0,x131})+$signed(-{1'b0,x67})+$signed(-{2'b0,x68}<<<3'd1)+$signed(-{1'b0,x292})+$signed(-{2'b0,x5}<<<3'd1)+$signed(-{1'b0,x357})+$signed(-{1'b0,x293})+$signed({3'b0,x166}<<<3'd2)+$signed({2'b0,x486}<<<3'd1)+$signed({1'b0,x294})+$signed({1'b0,x134})+$signed({3'b0,x359}<<<3'd2)+$signed({2'b0,x263}<<<3'd1)+$signed(-{1'b0,x358})+$signed(-{3'b0,x199}<<<3'd2)+$signed({3'b0,x424}<<<3'd2)+$signed(-{2'b0,x264}<<<3'd1)+$signed({1'b0,x8})+$signed({1'b0,x104})+$signed(-{1'b0,x328})+$signed(-{2'b0,x137}<<<3'd1)+$signed(-{2'b0,x235}<<<3'd1)+$signed({1'b0,x363})+$signed(-{1'b0,x427})+$signed({3'b0,x76}<<<3'd2)+$signed({1'b0,x300})+$signed({1'b0,x492})+$signed(-{1'b0,x460})+$signed({2'b0,x141}<<<3'd1)+$signed({2'b0,x493}<<<3'd1)+$signed({3'b0,x110}<<<3'd2)+$signed(-{1'b0,x462})+$signed({2'b0,x47}<<<3'd1)+$signed({3'b0,x177}<<<3'd2)+$signed({1'b0,x338})+$signed({2'b0,x467}<<<3'd1)+$signed(-{2'b0,x275}<<<3'd1)+$signed({2'b0,x372}<<<3'd1)+$signed({3'b0,x245}<<<3'd2)+$signed({2'b0,x213}<<<3'd1)+$signed({1'b0,x437})+$signed(-{2'b0,x181}<<<3'd1)+$signed(-{1'b0,x341})+$signed(-{3'b0,x438}<<<3'd2)+$signed(-{2'b0,x310}<<<3'd1)+$signed(-{2'b0,x470}<<<3'd1)+$signed({3'b0,x87}<<<3'd2)+$signed({2'b0,x407}<<<3'd1)+$signed({3'b0,x439}<<<3'd2)+$signed({2'b0,x471}<<<3'd1)+$signed({1'b0,x56})+$signed({3'b0,x377}<<<3'd2)+$signed({2'b0,x185}<<<3'd1)+$signed(-{1'b0,x89})+$signed({3'b0,x346}<<<3'd2)+$signed({3'b0,x378}<<<3'd2)+$signed({1'b0,x26})+$signed({1'b0,x122})+$signed({2'b0,x62}<<<3'd1)+$signed(-{2'b0,x315}<<<3'd1)+$signed({1'b0,x251})+$signed(-{2'b0,x27}<<<3'd1)+$signed({3'b0,x92}<<<3'd2)+$signed({3'b0,x95}<<<3'd2)+$signed(-{2'b0,x59}<<<3'd1)+$signed(-{2'b0,x379}<<<3'd1)+$signed({2'b0,x29}<<<3'd1)+$signed({2'b0,x125}<<<3'd1)+$signed({2'b0,x285}<<<3'd1)+$signed({3'b0,x94}<<<3'd2)+$signed({2'b0,x254}<<<3'd1)+$signed({3'b0,x415}<<<3'd2)+$signed({2'b0,x223}<<<3'd1);
assign sharing5 = $signed(-{3'b0,x192}<<<3'd2)+$signed({2'b0,x288}<<<3'd1)+$signed({2'b0,x290}<<<3'd1)+$signed({1'b0,x130})+$signed(-{1'b0,x162})+$signed(-{3'b0,x259}<<<3'd2)+$signed({3'b0,x422}<<<3'd2)+$signed({1'b0,x454})+$signed(-{2'b0,x423}<<<3'd1)+$signed({1'b0,x135})+$signed({3'b0,x265}<<<3'd2)+$signed({2'b0,x201}<<<3'd1)+$signed(-{3'b0,x457}<<<3'd2)+$signed(-{1'b0,x73})+$signed({3'b0,x394}<<<3'd2)+$signed(-{2'b0,x138}<<<3'd1)+$signed(-{2'b0,x447}<<<3'd1)+$signed(-{2'b0,x268}<<<3'd1)+$signed(-{3'b0,x174}<<<3'd2)+$signed({2'b0,x270}<<<3'd1)+$signed(-{1'b0,x302})+$signed(-{2'b0,x79}<<<3'd1)+$signed({1'b0,x463})+$signed({1'b0,x367})+$signed(-{3'b0,x464}<<<3'd2)+$signed(-{2'b0,x465}<<<3'd1)+$signed(-{1'b0,x337})+$signed({2'b0,x466}<<<3'd1)+$signed({3'b0,x435}<<<3'd2)+$signed({2'b0,x403}<<<3'd1)+$signed(-{3'b0,x84}<<<3'd2)+$signed(-{2'b0,x405}<<<3'd1)+$signed({1'b0,x53})+$signed({1'b0,x21})+$signed({1'b0,x149})+$signed({2'b0,x247}<<<3'd1)+$signed({2'b0,x279}<<<3'd1)+$signed(-{2'b0,x184}<<<3'd1)+$signed(-{2'b0,x345}<<<3'd1)+$signed({3'b0,x154}<<<3'd2)+$signed({3'b0,x220}<<<3'd2)+$signed({1'b0,x382})+$signed({3'b0,x191}<<<3'd2)+$signed({2'b0,x287}<<<3'd1);
assign sharing6 = $signed(-{3'b0,x448}<<<3'd2)+$signed({2'b0,x64}<<<3'd1)+$signed(-{1'b0,x320})+$signed(-{2'b0,x130}<<<3'd1)+$signed({1'b0,x195})+$signed(-{1'b0,x259})+$signed(-{3'b0,x68}<<<3'd2)+$signed(-{2'b0,x382}<<<3'd1)+$signed({3'b0,x70}<<<3'd2)+$signed(-{2'b0,x198}<<<3'd1)+$signed(-{1'b0,x454})+$signed(-{3'b0,x200}<<<3'd2)+$signed(-{1'b0,x136})+$signed({2'b0,x9}<<<3'd1)+$signed(-{2'b0,x202}<<<3'd1)+$signed(-{3'b0,x461}<<<3'd2)+$signed(-{2'b0,x333}<<<3'd1)+$signed({3'b0,x78}<<<3'd2)+$signed({2'b0,x79}<<<3'd1)+$signed(-{1'b0,x271})+$signed({1'b0,x16})+$signed(-{2'b0,x338}<<<3'd1)+$signed(-{4'b0,x403}<<<3'd3)+$signed(-{3'b0,x148}<<<3'd2)+$signed(-{1'b0,x468})+$signed(-{3'b0,x86}<<<3'd2)+$signed(-{1'b0,x22})+$signed({1'b0,x87})+$signed({2'b0,x24}<<<3'd1)+$signed(-{2'b0,x220}<<<3'd1)+$signed(-{3'b0,x30}<<<3'd2)+$signed({3'b0,x415}<<<3'd2)+$signed(-{3'b0,x288}<<<3'd2)+$signed(-{3'b0,x481}<<<3'd2)+$signed(-{3'b0,x417}<<<3'd2)+$signed({2'b0,x354}<<<3'd1)+$signed(-{4'b0,x165}<<<3'd3)+$signed(-{1'b0,x294})+$signed({2'b0,x423}<<<3'd1)+$signed(-{2'b0,x103}<<<3'd1)+$signed({3'b0,x424}<<<3'd2)+$signed({1'b0,x296})+$signed(-{3'b0,x233}<<<3'd2)+$signed({1'b0,x425})+$signed(-{2'b0,x235}<<<3'd1)+$signed({1'b0,x363})+$signed(-{3'b0,x494}<<<3'd2)+$signed(-{1'b0,x366})+$signed({3'b0,x432}<<<3'd2)+$signed(-{1'b0,x112})+$signed(-{3'b0,x305}<<<3'd2)+$signed(-{2'b0,x369}<<<3'd1)+$signed({2'b0,x114}<<<3'd1)+$signed(-{2'b0,x180}<<<3'd1)+$signed({1'b0,x372})+$signed({3'b0,x309}<<<3'd2)+$signed(-{2'b0,x53}<<<3'd1)+$signed({1'b0,x311})+$signed(-{3'b0,x184}<<<3'd2)+$signed(-{2'b0,x376}<<<3'd1)+$signed(-{3'b0,x442}<<<3'd2)+$signed({1'b0,x250})+$signed(-{3'b0,x379}<<<3'd2)+$signed(-{1'b0,x59})+$signed({2'b0,x254}<<<3'd1)+$signed(-{3'b0,x255}<<<3'd2);
assign sharing7 = $signed({3'b0,x192}<<<3'd2)+$signed({2'b0,x289}<<<3'd1)+$signed({2'b0,x385}<<<3'd1)+$signed({2'b0,x386}<<<3'd1)+$signed(-{2'b0,x2}<<<3'd1)+$signed(-{2'b0,x483}<<<3'd1)+$signed(-{2'b0,x3}<<<3'd1)+$signed(-{1'b0,x35})+$signed(-{2'b0,x228}<<<3'd1)+$signed({1'b0,x229})+$signed(-{3'b0,x422}<<<3'd2)+$signed(-{2'b0,x358}<<<3'd1)+$signed(-{3'b0,x39}<<<3'd2)+$signed({2'b0,x7}<<<3'd1)+$signed(-{1'b0,x359})+$signed(-{3'b0,x264}<<<3'd2)+$signed({2'b0,x328}<<<3'd1)+$signed({2'b0,x360}<<<3'd1)+$signed(-{2'b0,x104}<<<3'd1)+$signed(-{1'b0,x40})+$signed({1'b0,x105})+$signed({1'b0,x361})+$signed({1'b0,x394})+$signed(-{3'b0,x75}<<<3'd2)+$signed({1'b0,x428})+$signed(-{4'b0,x429}<<<3'd3)+$signed({2'b0,x302}<<<3'd1)+$signed(-{2'b0,x270}<<<3'd1)+$signed(-{1'b0,x206})+$signed({3'b0,x15}<<<3'd2)+$signed({3'b0,x399}<<<3'd2)+$signed({1'b0,x207})+$signed({1'b0,x175})+$signed(-{1'b0,x238})+$signed(-{3'b0,x304}<<<3'd2)+$signed(-{3'b0,x433}<<<3'd2)+$signed({2'b0,x178}<<<3'd1)+$signed(-{2'b0,x50}<<<3'd1)+$signed(-{3'b0,x115}<<<3'd2)+$signed(-{3'b0,x371}<<<3'd2)+$signed({1'b0,x339})+$signed({2'b0,x373}<<<3'd1)+$signed({3'b0,x151}<<<3'd2)+$signed(-{3'b0,x215}<<<3'd2)+$signed(-{2'b0,x247}<<<3'd1)+$signed(-{1'b0,x279})+$signed({2'b0,x248}<<<3'd1)+$signed(-{1'b0,x216})+$signed(-{3'b0,x57}<<<3'd2)+$signed({2'b0,x441}<<<3'd1)+$signed(-{3'b0,x281}<<<3'd2)+$signed(-{2'b0,x345}<<<3'd1)+$signed(-{2'b0,x314}<<<3'd1)+$signed(-{1'b0,x282})+$signed(-{2'b0,x346}<<<3'd1)+$signed({2'b0,x60}<<<3'd1)+$signed({2'b0,x125}<<<3'd1)+$signed({1'b0,x61})+$signed(-{2'b0,x286}<<<3'd1)+$signed(-{3'b0,x447}<<<3'd2);
assign sharing8 = $signed({3'b0,x160}<<<3'd2)+$signed(-{2'b0,x480}<<<3'd1)+$signed(-{3'b0,x353}<<<3'd2)+$signed({2'b0,x257}<<<3'd1)+$signed({1'b0,x1})+$signed({2'b0,x34}<<<3'd1)+$signed({2'b0,x130}<<<3'd1)+$signed(-{2'b0,x318}<<<3'd1)+$signed({2'b0,x485}<<<3'd1)+$signed(-{3'b0,x390}<<<3'd2)+$signed(-{3'b0,x230}<<<3'd2)+$signed(-{3'b0,x486}<<<3'd2)+$signed(-{3'b0,x167}<<<3'd2)+$signed(-{3'b0,x8}<<<3'd2)+$signed(-{3'b0,x72}<<<3'd2)+$signed({2'b0,x233}<<<3'd1)+$signed({4'b0,x43}<<<3'd3)+$signed({3'b0,x235}<<<3'd2)+$signed({2'b0,x75}<<<3'd1)+$signed({2'b0,x299}<<<3'd1)+$signed({3'b0,x331}<<<3'd2)+$signed(-{1'b0,x363})+$signed({1'b0,x76})+$signed({3'b0,x237}<<<3'd2)+$signed(-{2'b0,x13}<<<3'd1)+$signed({3'b0,x142}<<<3'd2)+$signed(-{3'b0,x206}<<<3'd2)+$signed(-{2'b0,x430}<<<3'd1)+$signed(-{3'b0,x431}<<<3'd2)+$signed(-{2'b0,x47}<<<3'd1)+$signed({1'b0,x143})+$signed(-{3'b0,x336}<<<3'd2)+$signed({3'b0,x370}<<<3'd2)+$signed(-{3'b0,x242}<<<3'd2)+$signed(-{3'b0,x466}<<<3'd2)+$signed(-{3'b0,x243}<<<3'd2)+$signed(-{2'b0,x211}<<<3'd1)+$signed({1'b0,x147})+$signed({3'b0,x212}<<<3'd2)+$signed(-{1'b0,x148})+$signed(-{1'b0,x437})+$signed({3'b0,x406}<<<3'd2)+$signed(-{1'b0,x61})+$signed({3'b0,x311}<<<3'd2)+$signed({3'b0,x312}<<<3'd2)+$signed({2'b0,x216}<<<3'd1)+$signed({2'b0,x190}<<<3'd1)+$signed(-{1'b0,x408})+$signed(-{3'b0,x474}<<<3'd2)+$signed(-{2'b0,x26}<<<3'd1)+$signed(-{1'b0,x154})+$signed(-{3'b0,x315}<<<3'd2)+$signed(-{2'b0,x411}<<<3'd1)+$signed({3'b0,x477}<<<3'd2)+$signed({2'b0,x349}<<<3'd1)+$signed(-{2'b0,x381}<<<3'd1)+$signed({2'b0,x446}<<<3'd1)+$signed(-{2'b0,x95}<<<3'd1);
assign sharing9 = $signed(-{1'b0,x320})+$signed({2'b0,x97}<<<3'd1)+$signed(-{2'b0,x449}<<<3'd1)+$signed(-{2'b0,x193}<<<3'd1)+$signed({3'b0,x226}<<<3'd2)+$signed(-{1'b0,x417})+$signed(-{2'b0,x2}<<<3'd1)+$signed(-{2'b0,x159}<<<3'd1)+$signed(-{3'b0,x355}<<<3'd2)+$signed(-{2'b0,x259}<<<3'd1)+$signed({1'b0,x227})+$signed(-{2'b0,x484}<<<3'd1)+$signed(-{1'b0,x36})+$signed(-{3'b0,x165}<<<3'd2)+$signed(-{3'b0,x38}<<<3'd2)+$signed(-{2'b0,x166}<<<3'd1)+$signed({4'b0,x455}<<<3'd3)+$signed({3'b0,x263}<<<3'd2)+$signed({3'b0,x71}<<<3'd2)+$signed(-{2'b0,x423}<<<3'd1)+$signed(-{2'b0,x359}<<<3'd1)+$signed({1'b0,x328})+$signed({3'b0,x137}<<<3'd2)+$signed({1'b0,x361})+$signed({3'b0,x395}<<<3'd2)+$signed(-{3'b0,x171}<<<3'd2)+$signed(-{3'b0,x44}<<<3'd2)+$signed(-{2'b0,x268}<<<3'd1)+$signed({1'b0,x332})+$signed({3'b0,x365}<<<3'd2)+$signed({2'b0,x461}<<<3'd1)+$signed(-{3'b0,x397}<<<3'd2)+$signed(-{2'b0,x301}<<<3'd1)+$signed({2'b0,x270}<<<3'd1)+$signed({2'b0,x78}<<<3'd1)+$signed(-{2'b0,x79}<<<3'd1)+$signed(-{2'b0,x207}<<<3'd1)+$signed(-{1'b0,x239})+$signed({3'b0,x400}<<<3'd2)+$signed({3'b0,x145}<<<3'd2)+$signed({1'b0,x177})+$signed({1'b0,x209})+$signed({2'b0,x51}<<<3'd1)+$signed({2'b0,x19}<<<3'd1)+$signed({1'b0,x115})+$signed({3'b0,x276}<<<3'd2)+$signed({2'b0,x244}<<<3'd1)+$signed({4'b0,x468}<<<3'd3)+$signed(-{2'b0,x307}<<<3'd1)+$signed(-{3'b0,x180}<<<3'd2)+$signed(-{3'b0,x469}<<<3'd2)+$signed({1'b0,x470})+$signed({3'b0,x55}<<<3'd2)+$signed({3'b0,x343}<<<3'd2)+$signed({1'b0,x151})+$signed(-{3'b0,x439}<<<3'd2)+$signed({3'b0,x280}<<<3'd2)+$signed(-{2'b0,x281}<<<3'd1)+$signed(-{1'b0,x441})+$signed({3'b0,x187}<<<3'd2)+$signed({2'b0,x27}<<<3'd1)+$signed(-{1'b0,x91})+$signed({3'b0,x380}<<<3'd2)+$signed(-{3'b0,x92}<<<3'd2)+$signed(-{3'b0,x157}<<<3'd2)+$signed(-{2'b0,x93}<<<3'd1)+$signed({2'b0,x223}<<<3'd1)+$signed({1'b0,x31});
assign sharing10 = $signed({3'b0,x128}<<<3'd2)+$signed(-{3'b0,x32}<<<3'd2)+$signed({3'b0,x289}<<<3'd2)+$signed({3'b0,x387}<<<3'd2)+$signed({2'b0,x483}<<<3'd1)+$signed({1'b0,x419})+$signed(-{3'b0,x323}<<<3'd2)+$signed({3'b0,x484}<<<3'd2)+$signed(-{1'b0,x451})+$signed(-{3'b0,x420}<<<3'd2)+$signed(-{1'b0,x260})+$signed({2'b0,x197}<<<3'd1)+$signed(-{2'b0,x293}<<<3'd1)+$signed(-{4'b0,x134}<<<3'd3)+$signed(-{1'b0,x422})+$signed({2'b0,x423}<<<3'd1)+$signed(-{1'b0,x7})+$signed({1'b0,x488})+$signed({3'b0,x393}<<<3'd2)+$signed(-{3'b0,x73}<<<3'd2)+$signed(-{1'b0,x233})+$signed({3'b0,x490}<<<3'd2)+$signed(-{1'b0,x426})+$signed({3'b0,x43}<<<3'd2)+$signed({3'b0,x235}<<<3'd2)+$signed(-{3'b0,x171}<<<3'd2)+$signed(-{4'b0,x44}<<<3'd3)+$signed({3'b0,x364}<<<3'd2)+$signed({3'b0,x460}<<<3'd2)+$signed(-{2'b0,x140}<<<3'd1)+$signed({2'b0,x269}<<<3'd1)+$signed(-{3'b0,x366}<<<3'd2)+$signed({2'b0,x78}<<<3'd1)+$signed({3'b0,x79}<<<3'd2)+$signed({3'b0,x208}<<<3'd2)+$signed(-{3'b0,x18}<<<3'd2)+$signed({2'b0,x178}<<<3'd1)+$signed({1'b0,x210})+$signed(-{3'b0,x306}<<<3'd2)+$signed({3'b0,x115}<<<3'd2)+$signed(-{3'b0,x402}<<<3'd2)+$signed(-{3'b0,x51}<<<3'd2)+$signed({3'b0,x468}<<<3'd2)+$signed({3'b0,x245}<<<3'd2)+$signed(-{1'b0,x213})+$signed({2'b0,x406}<<<3'd1)+$signed(-{1'b0,x182})+$signed(-{4'b0,x279}<<<3'd3)+$signed(-{2'b0,x247}<<<3'd1)+$signed(-{3'b0,x440}<<<3'd2)+$signed({2'b0,x24}<<<3'd1)+$signed({1'b0,x88})+$signed({2'b0,x216}<<<3'd1)+$signed(-{2'b0,x152}<<<3'd1)+$signed(-{1'b0,x376})+$signed({1'b0,x57})+$signed(-{3'b0,x153}<<<3'd2)+$signed(-{2'b0,x217}<<<3'd1)+$signed({2'b0,x410}<<<3'd1)+$signed(-{2'b0,x91}<<<3'd1)+$signed({3'b0,x124}<<<3'd2)+$signed({3'b0,x158}<<<3'd2)+$signed(-{1'b0,x60})+$signed({3'b0,x93}<<<3'd2)+$signed({2'b0,x477}<<<3'd1)+$signed(-{4'b0,x62}<<<3'd3)+$signed({3'b0,x126}<<<3'd2)+$signed({2'b0,x254}<<<3'd1)+$signed({3'b0,x191}<<<3'd2)+$signed(-{2'b0,x319}<<<3'd1);
assign sharing11 = $signed(-{3'b0,x480}<<<3'd2)+$signed(-{3'b0,x161}<<<3'd2)+$signed({3'b0,x66}<<<3'd2)+$signed({3'b0,x162}<<<3'd2)+$signed(-{3'b0,x98}<<<3'd2)+$signed(-{2'b0,x226}<<<3'd1)+$signed({2'b0,x67}<<<3'd1)+$signed({1'b0,x259})+$signed({1'b0,x131})+$signed({2'b0,x228}<<<3'd1)+$signed(-{2'b0,x196}<<<3'd1)+$signed({2'b0,x485}<<<3'd1)+$signed(-{2'b0,x358}<<<3'd1)+$signed(-{1'b0,x6})+$signed(-{3'b0,x295}<<<3'd2)+$signed({2'b0,x391}<<<3'd1)+$signed(-{1'b0,x168})+$signed(-{1'b0,x424})+$signed({2'b0,x361}<<<3'd1)+$signed(-{2'b0,x105}<<<3'd1)+$signed(-{1'b0,x169})+$signed(-{1'b0,x74})+$signed(-{2'b0,x139}<<<3'd1)+$signed(-{2'b0,x447}<<<3'd1)+$signed({3'b0,x76}<<<3'd2)+$signed({2'b0,x268}<<<3'd1)+$signed(-{3'b0,x46}<<<3'd2)+$signed({2'b0,x302}<<<3'd1)+$signed({2'b0,x398}<<<3'd1)+$signed({4'b0,x495}<<<3'd3)+$signed(-{1'b0,x206})+$signed(-{2'b0,x431}<<<3'd1)+$signed(-{1'b0,x368})+$signed({3'b0,x274}<<<3'd2)+$signed(-{2'b0,x466}<<<3'd1)+$signed(-{2'b0,x179}<<<3'd1)+$signed({3'b0,x20}<<<3'd2)+$signed(-{3'b0,x118}<<<3'd2)+$signed(-{2'b0,x438}<<<3'd1)+$signed({3'b0,x407}<<<3'd2)+$signed({2'b0,x151}<<<3'd1)+$signed(-{1'b0,x56})+$signed(-{3'b0,x345}<<<3'd2)+$signed(-{1'b0,x249})+$signed(-{2'b0,x218}<<<3'd1)+$signed(-{2'b0,x346}<<<3'd1)+$signed({3'b0,x443}<<<3'd2)+$signed({2'b0,x59}<<<3'd1)+$signed({1'b0,x27})+$signed({2'b0,x123}<<<3'd1)+$signed(-{3'b0,x28}<<<3'd2)+$signed(-{3'b0,x156}<<<3'd2)+$signed(-{1'b0,x380})+$signed(-{3'b0,x125}<<<3'd2)+$signed({2'b0,x61}<<<3'd1)+$signed({1'b0,x445})+$signed({3'b0,x446}<<<3'd2)+$signed({2'b0,x222}<<<3'd1)+$signed(-{2'b0,x415}<<<3'd1);
assign sharing12 = $signed({3'b0,x384}<<<3'd2)+$signed({2'b0,x288}<<<3'd1)+$signed(-{2'b0,x256}<<<3'd1)+$signed({3'b0,x481}<<<3'd2)+$signed({3'b0,x418}<<<3'd2)+$signed(-{3'b0,x99}<<<3'd2)+$signed({2'b0,x419}<<<3'd1)+$signed(-{2'b0,x195}<<<3'd1)+$signed(-{2'b0,x3}<<<3'd1)+$signed({3'b0,x292}<<<3'd2)+$signed({3'b0,x420}<<<3'd2)+$signed(-{1'b0,x35})+$signed(-{2'b0,x227}<<<3'd1)+$signed({3'b0,x37}<<<3'd2)+$signed(-{3'b0,x261}<<<3'd2)+$signed({3'b0,x70}<<<3'd2)+$signed({2'b0,x390}<<<3'd1)+$signed({3'b0,x262}<<<3'd2)+$signed(-{2'b0,x166}<<<3'd1)+$signed(-{2'b0,x287}<<<3'd1)+$signed({2'b0,x167}<<<3'd1)+$signed({2'b0,x423}<<<3'd1)+$signed({2'b0,x327}<<<3'd1)+$signed(-{2'b0,x487}<<<3'd1)+$signed({2'b0,x296}<<<3'd1)+$signed({2'b0,x456}<<<3'd1)+$signed(-{1'b0,x328})+$signed({3'b0,x361}<<<3'd2)+$signed({2'b0,x73}<<<3'd1)+$signed({2'b0,x297}<<<3'd1)+$signed(-{1'b0,x169})+$signed({2'b0,x202}<<<3'd1)+$signed({2'b0,x426}<<<3'd1)+$signed(-{1'b0,x298})+$signed({3'b0,x75}<<<3'd2)+$signed({1'b0,x43})+$signed({1'b0,x427})+$signed({3'b0,x364}<<<3'd2)+$signed(-{2'b0,x428}<<<3'd1)+$signed(-{3'b0,x45}<<<3'd2)+$signed(-{2'b0,x269}<<<3'd1)+$signed({3'b0,x78}<<<3'd2)+$signed({3'b0,x15}<<<3'd2)+$signed(-{2'b0,x239}<<<3'd1)+$signed(-{3'b0,x144}<<<3'd2)+$signed({2'b0,x400}<<<3'd1)+$signed({1'b0,x432})+$signed({3'b0,x145}<<<3'd2)+$signed({3'b0,x402}<<<3'd2)+$signed({1'b0,x146})+$signed({1'b0,x274})+$signed({3'b0,x19}<<<3'd2)+$signed(-{2'b0,x403}<<<3'd1)+$signed(-{2'b0,x372}<<<3'd1)+$signed(-{1'b0,x20})+$signed(-{1'b0,x308})+$signed({3'b0,x55}<<<3'd2)+$signed({3'b0,x407}<<<3'd2)+$signed({3'b0,x439}<<<3'd2)+$signed(-{2'b0,x184}<<<3'd1)+$signed(-{2'b0,x344}<<<3'd1)+$signed({3'b0,x345}<<<3'd2)+$signed({2'b0,x121}<<<3'd1)+$signed({2'b0,x185}<<<3'd1)+$signed(-{3'b0,x313}<<<3'd2)+$signed(-{3'b0,x474}<<<3'd2)+$signed({2'b0,x58}<<<3'd1)+$signed(-{1'b0,x250})+$signed({2'b0,x91}<<<3'd1)+$signed({2'b0,x219}<<<3'd1)+$signed({2'b0,x347}<<<3'd1)+$signed({3'b0,x156}<<<3'd2)+$signed({3'b0,x316}<<<3'd2)+$signed(-{2'b0,x59}<<<3'd1)+$signed(-{1'b0,x411})+$signed(-{3'b0,x252}<<<3'd2)+$signed(-{2'b0,x124}<<<3'd1)+$signed(-{3'b0,x478}<<<3'd2)+$signed({2'b0,x127}<<<3'd1)+$signed(-{1'b0,x319});
assign sharing13 = $signed({2'b0,x0}<<<3'd1)+$signed({2'b0,x320}<<<3'd1)+$signed({2'b0,x224}<<<3'd1)+$signed(-{1'b0,x128})+$signed({2'b0,x321}<<<3'd1)+$signed(-{2'b0,x193}<<<3'd1)+$signed(-{3'b0,x98}<<<3'd2)+$signed(-{3'b0,x163}<<<3'd2)+$signed({2'b0,x36}<<<3'd1)+$signed({1'b0,x132})+$signed(-{3'b0,x358}<<<3'd2)+$signed({1'b0,x455})+$signed(-{3'b0,x457}<<<3'd2)+$signed(-{3'b0,x395}<<<3'd2)+$signed({2'b0,x492}<<<3'd1)+$signed(-{2'b0,x396}<<<3'd1)+$signed(-{2'b0,x109}<<<3'd1)+$signed(-{3'b0,x430}<<<3'd2)+$signed({2'b0,x463}<<<3'd1)+$signed(-{2'b0,x303}<<<3'd1)+$signed({2'b0,x336}<<<3'd1)+$signed({2'b0,x49}<<<3'd1)+$signed({1'b0,x177})+$signed({2'b0,x401}<<<3'd1)+$signed({3'b0,x114}<<<3'd2)+$signed({2'b0,x306}<<<3'd1)+$signed({2'b0,x433}<<<3'd1)+$signed(-{1'b0,x369})+$signed(-{3'b0,x210}<<<3'd2)+$signed({2'b0,x467}<<<3'd1)+$signed(-{3'b0,x370}<<<3'd2)+$signed(-{1'b0,x373})+$signed(-{1'b0,x277})+$signed({2'b0,x278}<<<3'd1)+$signed(-{2'b0,x119}<<<3'd1)+$signed(-{1'b0,x87})+$signed(-{2'b0,x280}<<<3'd1)+$signed(-{2'b0,x312}<<<3'd1)+$signed(-{2'b0,x377}<<<3'd1)+$signed(-{1'b0,x158})+$signed({2'b0,x315}<<<3'd1)+$signed(-{1'b0,x123})+$signed({2'b0,x476}<<<3'd1)+$signed(-{2'b0,x189}<<<3'd1)+$signed(-{1'b0,x253})+$signed({3'b0,x382}<<<3'd2)+$signed(-{2'b0,x446}<<<3'd1)+$signed({1'b0,x126})+$signed({3'b0,x95}<<<3'd2)+$signed({2'b0,x31}<<<3'd1)+$signed({1'b0,x383});
assign sharing14 = $signed({3'b0,x416}<<<3'd2)+$signed(-{3'b0,x256}<<<3'd2)+$signed({2'b0,x289}<<<3'd1)+$signed({1'b0,x130})+$signed({3'b0,x483}<<<3'd2)+$signed({2'b0,x163}<<<3'd1)+$signed({2'b0,x387}<<<3'd1)+$signed({3'b0,x196}<<<3'd2)+$signed({2'b0,x164}<<<3'd1)+$signed({1'b0,x68})+$signed(-{2'b0,x389}<<<3'd1)+$signed(-{3'b0,x486}<<<3'd2)+$signed({2'b0,x358}<<<3'd1)+$signed(-{1'b0,x38})+$signed({3'b0,x455}<<<3'd2)+$signed({3'b0,x263}<<<3'd2)+$signed({3'b0,x295}<<<3'd2)+$signed({3'b0,x167}<<<3'd2)+$signed({3'b0,x136}<<<3'd2)+$signed({3'b0,x296}<<<3'd2)+$signed({1'b0,x72})+$signed(-{3'b0,x487}<<<3'd2)+$signed({3'b0,x415}<<<3'd2)+$signed(-{1'b0,x359})+$signed(-{3'b0,x137}<<<3'd2)+$signed(-{1'b0,x425})+$signed({3'b0,x266}<<<3'd2)+$signed(-{1'b0,x490})+$signed({3'b0,x331}<<<3'd2)+$signed({2'b0,x139}<<<3'd1)+$signed(-{3'b0,x75}<<<3'd2)+$signed({3'b0,x492}<<<3'd2)+$signed(-{3'b0,x12}<<<3'd2)+$signed(-{1'b0,x268})+$signed({3'b0,x205}<<<3'd2)+$signed(-{2'b0,x13}<<<3'd1)+$signed(-{1'b0,x45})+$signed({3'b0,x270}<<<3'd2)+$signed({2'b0,x46}<<<3'd1)+$signed({2'b0,x334}<<<3'd1)+$signed({2'b0,x462}<<<3'd1)+$signed(-{2'b0,x494}<<<3'd1)+$signed(-{2'b0,x14}<<<3'd1)+$signed(-{2'b0,x302}<<<3'd1)+$signed(-{2'b0,x176}<<<3'd1)+$signed({2'b0,x241}<<<3'd1)+$signed({3'b0,x50}<<<3'd2)+$signed(-{2'b0,x210}<<<3'd1)+$signed({2'b0,x83}<<<3'd1)+$signed({2'b0,x148}<<<3'd1)+$signed(-{2'b0,x84}<<<3'd1)+$signed(-{3'b0,x21}<<<3'd2)+$signed({2'b0,x373}<<<3'd1)+$signed({3'b0,x470}<<<3'd2)+$signed(-{2'b0,x342}<<<3'd1)+$signed({1'b0,x246})+$signed({3'b0,x248}<<<3'd2)+$signed({2'b0,x152}<<<3'd1)+$signed({3'b0,x281}<<<3'd2)+$signed(-{2'b0,x377}<<<3'd1)+$signed(-{2'b0,x282}<<<3'd1)+$signed({1'b0,x218})+$signed(-{2'b0,x474}<<<3'd1)+$signed({3'b0,x443}<<<3'd2)+$signed({2'b0,x475}<<<3'd1)+$signed(-{1'b0,x27})+$signed(-{1'b0,x445})+$signed(-{1'b0,x478})+$signed({3'b0,x447}<<<3'd2)+$signed(-{2'b0,x127}<<<3'd1);
assign sharing15 = $signed(-{2'b0,x448}<<<3'd1)+$signed(-{2'b0,x128}<<<3'd1)+$signed(-{1'b0,x384})+$signed({3'b0,x449}<<<3'd2)+$signed({2'b0,x193}<<<3'd1)+$signed(-{1'b0,x65})+$signed(-{1'b0,x381})+$signed({2'b0,x322}<<<3'd1)+$signed({2'b0,x323}<<<3'd1)+$signed(-{1'b0,x451})+$signed(-{3'b0,x69}<<<3'd2)+$signed(-{3'b0,x197}<<<3'd2)+$signed(-{2'b0,x255}<<<3'd1)+$signed({1'b0,x198})+$signed(-{1'b0,x70})+$signed({3'b0,x392}<<<3'd2)+$signed(-{2'b0,x200}<<<3'd1)+$signed(-{2'b0,x265}<<<3'd1)+$signed(-{3'b0,x267}<<<3'd2)+$signed({2'b0,x396}<<<3'd1)+$signed({1'b0,x204})+$signed(-{3'b0,x141}<<<3'd2)+$signed(-{2'b0,x461}<<<3'd1)+$signed(-{2'b0,x206}<<<3'd1)+$signed(-{3'b0,x335}<<<3'd2)+$signed(-{3'b0,x336}<<<3'd2)+$signed({2'b0,x272}<<<3'd1)+$signed(-{2'b0,x80}<<<3'd1)+$signed(-{2'b0,x402}<<<3'd1)+$signed(-{3'b0,x468}<<<3'd2)+$signed(-{2'b0,x340}<<<3'd1)+$signed(-{1'b0,x404})+$signed(-{2'b0,x473}<<<3'd1)+$signed({1'b0,x345})+$signed({1'b0,x409})+$signed(-{2'b0,x346}<<<3'd1)+$signed({1'b0,x283})+$signed({2'b0,x157}<<<3'd1)+$signed({2'b0,x285}<<<3'd1)+$signed(-{2'b0,x477}<<<3'd1)+$signed(-{1'b0,x350})+$signed(-{2'b0,x33}<<<3'd1)+$signed(-{2'b0,x353}<<<3'd1)+$signed(-{3'b0,x226}<<<3'd2)+$signed({2'b0,x355}<<<3'd1)+$signed({3'b0,x229}<<<3'd2)+$signed({3'b0,x357}<<<3'd2)+$signed({2'b0,x421}<<<3'd1)+$signed(-{1'b0,x298})+$signed({3'b0,x427}<<<3'd2)+$signed({3'b0,x493}<<<3'd2)+$signed(-{3'b0,x111}<<<3'd2)+$signed(-{1'b0,x113})+$signed({2'b0,x242}<<<3'd1)+$signed(-{2'b0,x114}<<<3'd1)+$signed({2'b0,x180}<<<3'd1)+$signed(-{1'b0,x372})+$signed(-{3'b0,x118}<<<3'd2)+$signed(-{3'b0,x439}<<<3'd2)+$signed({2'b0,x119}<<<3'd1)+$signed(-{3'b0,x184}<<<3'd2)+$signed({2'b0,x312}<<<3'd1)+$signed({3'b0,x188}<<<3'd2)+$signed(-{1'b0,x125})+$signed({2'b0,x63}<<<3'd1);
assign sharing16 = $signed({2'b0,x256}<<<3'd1)+$signed({2'b0,x65}<<<3'd1)+$signed({2'b0,x385}<<<3'd1)+$signed(-{2'b0,x449}<<<3'd1)+$signed({2'b0,x451}<<<3'd1)+$signed(-{2'b0,x131}<<<3'd1)+$signed({2'b0,x68}<<<3'd1)+$signed(-{2'b0,x388}<<<3'd1)+$signed({2'b0,x389}<<<3'd1)+$signed(-{2'b0,x133}<<<3'd1)+$signed(-{1'b0,x325})+$signed({3'b0,x390}<<<3'd2)+$signed(-{1'b0,x454})+$signed({3'b0,x391}<<<3'd2)+$signed({2'b0,x71}<<<3'd1)+$signed(-{2'b0,x455}<<<3'd1)+$signed(-{2'b0,x72}<<<3'd1)+$signed(-{2'b0,x392}<<<3'd1)+$signed(-{2'b0,x9}<<<3'd1)+$signed({3'b0,x75}<<<3'd2)+$signed(-{2'b0,x139}<<<3'd1)+$signed({3'b0,x76}<<<3'd2)+$signed(-{2'b0,x332}<<<3'd1)+$signed({2'b0,x141}<<<3'd1)+$signed({2'b0,x269}<<<3'd1)+$signed(-{2'b0,x205}<<<3'd1)+$signed({2'b0,x142}<<<3'd1)+$signed(-{2'b0,x398}<<<3'd1)+$signed(-{2'b0,x207}<<<3'd1)+$signed({2'b0,x17}<<<3'd1)+$signed({2'b0,x209}<<<3'd1)+$signed(-{1'b0,x82})+$signed(-{3'b0,x275}<<<3'd2)+$signed({3'b0,x212}<<<3'd2)+$signed({2'b0,x21}<<<3'd1)+$signed({1'b0,x213})+$signed(-{2'b0,x150}<<<3'd1)+$signed(-{2'b0,x406}<<<3'd1)+$signed({3'b0,x215}<<<3'd2)+$signed({2'b0,x151}<<<3'd1)+$signed(-{2'b0,x279}<<<3'd1)+$signed(-{1'b0,x24})+$signed(-{1'b0,x88})+$signed({2'b0,x282}<<<3'd1)+$signed({2'b0,x346}<<<3'd1)+$signed(-{2'b0,x283}<<<3'd1)+$signed(-{2'b0,x411}<<<3'd1)+$signed({2'b0,x220}<<<3'd1)+$signed({1'b0,x476})+$signed({2'b0,x93}<<<3'd1)+$signed({1'b0,x29})+$signed({3'b0,x30}<<<3'd2)+$signed({1'b0,x352})+$signed(-{1'b0,x225})+$signed(-{3'b0,x162}<<<3'd2)+$signed(-{1'b0,x34})+$signed({3'b0,x292}<<<3'd2)+$signed({3'b0,x484}<<<3'd2)+$signed({1'b0,x228})+$signed(-{2'b0,x37}<<<3'd1)+$signed(-{2'b0,x422}<<<3'd1)+$signed({1'b0,x361})+$signed({1'b0,x489})+$signed({3'b0,x362}<<<3'd2)+$signed(-{2'b0,x236}<<<3'd1)+$signed(-{1'b0,x108})+$signed(-{3'b0,x45}<<<3'd2)+$signed(-{2'b0,x493}<<<3'd1)+$signed({3'b0,x238}<<<3'd2)+$signed({2'b0,x111}<<<3'd1)+$signed({2'b0,x431}<<<3'd1)+$signed({4'b0,x112}<<<3'd3)+$signed({3'b0,x176}<<<3'd2)+$signed({2'b0,x305}<<<3'd1)+$signed({2'b0,x114}<<<3'd1)+$signed(-{2'b0,x244}<<<3'd1)+$signed(-{2'b0,x436}<<<3'd1)+$signed(-{3'b0,x118}<<<3'd2)+$signed({2'b0,x54}<<<3'd1)+$signed(-{1'b0,x248})+$signed({3'b0,x58}<<<3'd2)+$signed({2'b0,x378}<<<3'd1)+$signed(-{2'b0,x442}<<<3'd1)+$signed({3'b0,x443}<<<3'd2)+$signed({3'b0,x316}<<<3'd2)+$signed({4'b0,x381}<<<3'd3)+$signed({2'b0,x63}<<<3'd1);
assign sharing17 = $signed({3'b0,x448}<<<3'd2)+$signed({2'b0,x96}<<<3'd1)+$signed(-{3'b0,x193}<<<3'd2)+$signed({3'b0,x98}<<<3'd2)+$signed({1'b0,x482})+$signed(-{1'b0,x67})+$signed({2'b0,x260}<<<3'd1)+$signed({1'b0,x420})+$signed(-{2'b0,x4}<<<3'd1)+$signed({3'b0,x69}<<<3'd2)+$signed(-{2'b0,x421}<<<3'd1)+$signed(-{3'b0,x102}<<<3'd2)+$signed({2'b0,x294}<<<3'd1)+$signed({3'b0,x7}<<<3'd2)+$signed(-{2'b0,x103}<<<3'd1)+$signed({3'b0,x104}<<<3'd2)+$signed({1'b0,x488})+$signed(-{2'b0,x105}<<<3'd1)+$signed(-{1'b0,x41})+$signed(-{1'b0,x457})+$signed({1'b0,x234})+$signed(-{1'b0,x10})+$signed(-{1'b0,x266})+$signed({2'b0,x427}<<<3'd1)+$signed(-{3'b0,x331}<<<3'd2)+$signed(-{2'b0,x363}<<<3'd1)+$signed(-{2'b0,x300}<<<3'd1)+$signed({2'b0,x77}<<<3'd1)+$signed({2'b0,x333}<<<3'd1)+$signed(-{2'b0,x237}<<<3'd1)+$signed({2'b0,x14}<<<3'd1)+$signed(-{3'b0,x175}<<<3'd2)+$signed(-{1'b0,x239})+$signed({2'b0,x145}<<<3'd1)+$signed(-{1'b0,x148})+$signed({1'b0,x181})+$signed(-{1'b0,x437})+$signed(-{2'b0,x182}<<<3'd1)+$signed(-{2'b0,x214}<<<3'd1)+$signed(-{2'b0,x86}<<<3'd1)+$signed(-{2'b0,x87}<<<3'd1)+$signed(-{2'b0,x55}<<<3'd1)+$signed({2'b0,x56}<<<3'd1)+$signed({1'b0,x152})+$signed({2'b0,x475}<<<3'd1)+$signed({3'b0,x28}<<<3'd2)+$signed(-{2'b0,x126}<<<3'd1)+$signed(-{1'b0,x284})+$signed(-{1'b0,x380})+$signed(-{3'b0,x317}<<<3'd2)+$signed({2'b0,x286}<<<3'd1);
assign sharing18 = $signed({3'b0,x224}<<<3'd2)+$signed({2'b0,x385}<<<3'd1)+$signed(-{2'b0,x417}<<<3'd1)+$signed({3'b0,x418}<<<3'd2)+$signed({2'b0,x290}<<<3'd1)+$signed({1'b0,x34})+$signed({1'b0,x130})+$signed({3'b0,x131}<<<3'd2)+$signed({1'b0,x258})+$signed(-{1'b0,x35})+$signed({3'b0,x164}<<<3'd2)+$signed({3'b0,x356}<<<3'd2)+$signed(-{1'b0,x228})+$signed({3'b0,x229}<<<3'd2)+$signed({2'b0,x421}<<<3'd1)+$signed({3'b0,x358}<<<3'd2)+$signed({3'b0,x102}<<<3'd2)+$signed({1'b0,x166})+$signed(-{3'b0,x231}<<<3'd2)+$signed({2'b0,x199}<<<3'd1)+$signed({2'b0,x360}<<<3'd1)+$signed({1'b0,x232})+$signed({2'b0,x106}<<<3'd1)+$signed({3'b0,x267}<<<3'd2)+$signed(-{1'b0,x11})+$signed({3'b0,x172}<<<3'd2)+$signed({2'b0,x492}<<<3'd1)+$signed(-{1'b0,x460})+$signed({3'b0,x109}<<<3'd2)+$signed({1'b0,x141})+$signed({2'b0,x302}<<<3'd1)+$signed({1'b0,x366})+$signed({2'b0,x430}<<<3'd1)+$signed({3'b0,x463}<<<3'd2)+$signed(-{3'b0,x111}<<<3'd2)+$signed(-{2'b0,x79}<<<3'd1)+$signed(-{1'b0,x367})+$signed({2'b0,x16}<<<3'd1)+$signed({2'b0,x80}<<<3'd1)+$signed({1'b0,x368})+$signed({2'b0,x432}<<<3'd1)+$signed({2'b0,x273}<<<3'd1)+$signed(-{1'b0,x272})+$signed(-{3'b0,x274}<<<3'd2)+$signed({2'b0,x51}<<<3'd1)+$signed(-{2'b0,x339}<<<3'd1)+$signed({3'b0,x276}<<<3'd2)+$signed({2'b0,x372}<<<3'd1)+$signed(-{3'b0,x404}<<<3'd2)+$signed(-{2'b0,x117}<<<3'd1)+$signed({3'b0,x278}<<<3'd2)+$signed({2'b0,x374}<<<3'd1)+$signed({3'b0,x406}<<<3'd2)+$signed(-{2'b0,x246}<<<3'd1)+$signed(-{1'b0,x310})+$signed({2'b0,x55}<<<3'd1)+$signed({1'b0,x87})+$signed({1'b0,x183})+$signed({3'b0,x152}<<<3'd2)+$signed({4'b0,x408}<<<3'd3)+$signed({1'b0,x88})+$signed({2'b0,x440}<<<3'd1)+$signed({3'b0,x472}<<<3'd2)+$signed(-{2'b0,x439}<<<3'd1)+$signed({1'b0,x409})+$signed({3'b0,x378}<<<3'd2)+$signed(-{2'b0,x26}<<<3'd1)+$signed({1'b0,x282})+$signed({3'b0,x91}<<<3'd2)+$signed({1'b0,x221})+$signed(-{1'b0,x59})+$signed(-{3'b0,x220}<<<3'd2)+$signed({2'b0,x284}<<<3'd1)+$signed({1'b0,x316})+$signed({2'b0,x412}<<<3'd1)+$signed({3'b0,x317}<<<3'd2)+$signed({2'b0,x381}<<<3'd1)+$signed({1'b0,x253})+$signed(-{2'b0,x445}<<<3'd1)+$signed({3'b0,x222}<<<3'd2)+$signed({1'b0,x62})+$signed({2'b0,x255}<<<3'd1);
assign sharing19 = $signed(-{3'b0,x192}<<<3'd2)+$signed({2'b0,x129}<<<3'd1)+$signed(-{2'b0,x481}<<<3'd1)+$signed(-{2'b0,x482}<<<3'd1)+$signed({1'b0,x450})+$signed(-{3'b0,x483}<<<3'd2)+$signed(-{2'b0,x484}<<<3'd1)+$signed({1'b0,x350})+$signed({3'b0,x197}<<<3'd2)+$signed({2'b0,x389}<<<3'd1)+$signed(-{3'b0,x325}<<<3'd2)+$signed(-{2'b0,x70}<<<3'd1)+$signed({1'b0,x486})+$signed({1'b0,x134})+$signed(-{2'b0,x294}<<<3'd1)+$signed({2'b0,x167}<<<3'd1)+$signed({3'b0,x136}<<<3'd2)+$signed({2'b0,x392}<<<3'd1)+$signed(-{1'b0,x488})+$signed({2'b0,x73}<<<3'd1)+$signed(-{2'b0,x425}<<<3'd1)+$signed(-{3'b0,x138}<<<3'd2)+$signed({1'b0,x74})+$signed(-{1'b0,x170})+$signed(-{1'b0,x298})+$signed({2'b0,x269}<<<3'd1)+$signed({1'b0,x77})+$signed({2'b0,x110}<<<3'd1)+$signed({2'b0,x46}<<<3'd1)+$signed(-{2'b0,x142}<<<3'd1)+$signed(-{2'b0,x174}<<<3'd1)+$signed({2'b0,x335}<<<3'd1)+$signed(-{3'b0,x399}<<<3'd2)+$signed(-{2'b0,x47}<<<3'd1)+$signed({2'b0,x208}<<<3'd1)+$signed({1'b0,x144})+$signed(-{2'b0,x400}<<<3'd1)+$signed(-{2'b0,x464}<<<3'd1)+$signed({2'b0,x145}<<<3'd1)+$signed({1'b0,x177})+$signed({3'b0,x82}<<<3'd2)+$signed(-{2'b0,x306}<<<3'd1)+$signed(-{2'b0,x148}<<<3'd1)+$signed({1'b0,x212})+$signed({1'b0,x308})+$signed(-{1'b0,x436})+$signed(-{2'b0,x438}<<<3'd1)+$signed(-{1'b0,x86})+$signed(-{3'b0,x30}<<<3'd2)+$signed({3'b0,x217}<<<3'd2)+$signed({2'b0,x185}<<<3'd1)+$signed(-{1'b0,x473})+$signed({3'b0,x154}<<<3'd2)+$signed(-{3'b0,x90}<<<3'd2)+$signed({2'b0,x251}<<<3'd1)+$signed(-{1'b0,x283})+$signed(-{3'b0,x380}<<<3'd2)+$signed(-{3'b0,x190}<<<3'd2)+$signed(-{2'b0,x158}<<<3'd1)+$signed({1'b0,x478})+$signed(-{2'b0,x223}<<<3'd1);
assign sharing20 = $signed(-{2'b0,x464}<<<3'd1)+$signed(-{1'b0,x257})+$signed({1'b0,x34})+$signed(-{1'b0,x290})+$signed({1'b0,x275})+$signed(-{3'b0,x5}<<<3'd2)+$signed({2'b0,x437}<<<3'd1)+$signed({1'b0,x405})+$signed(-{3'b0,x230}<<<3'd2)+$signed(-{2'b0,x215}<<<3'd1)+$signed({3'b0,x8}<<<3'd2)+$signed({3'b0,x168}<<<3'd2)+$signed(-{1'b0,x24})+$signed(-{1'b0,x57})+$signed(-{1'b0,x217})+$signed({3'b0,x330}<<<3'd2)+$signed(-{2'b0,x378}<<<3'd1)+$signed(-{1'b0,x410})+$signed(-{3'b0,x491}<<<3'd2)+$signed({2'b0,x44}<<<3'd1)+$signed(-{2'b0,x140}<<<3'd1)+$signed(-{2'b0,x220}<<<3'd1)+$signed({3'b0,x61}<<<3'd2)+$signed(-{4'b0,x286}<<<3'd3)+$signed({3'b0,x62}<<<3'd2)+$signed({1'b0,x30})+$signed(-{2'b0,x143}<<<3'd1);
assign sharing21 = $signed(-{3'b0,x81}<<<3'd2)+$signed({2'b0,x161}<<<3'd1)+$signed(-{3'b0,x159}<<<3'd2)+$signed({1'b0,x338})+$signed(-{3'b0,x179}<<<3'd2)+$signed({2'b0,x147}<<<3'd1)+$signed({1'b0,x291})+$signed({2'b0,x67}<<<3'd1)+$signed(-{3'b0,x259}<<<3'd2)+$signed(-{1'b0,x243})+$signed(-{3'b0,x100}<<<3'd2)+$signed(-{2'b0,x452}<<<3'd1)+$signed(-{3'b0,x214}<<<3'd2)+$signed({2'b0,x86}<<<3'd1)+$signed(-{3'b0,x135}<<<3'd2)+$signed(-{3'b0,x247}<<<3'd2)+$signed(-{1'b0,x311})+$signed(-{2'b0,x40}<<<3'd1)+$signed({1'b0,x216})+$signed(-{1'b0,x376})+$signed(-{3'b0,x153}<<<3'd2)+$signed(-{2'b0,x41}<<<3'd1)+$signed({1'b0,x233})+$signed(-{3'b0,x25}<<<3'd2)+$signed({3'b0,x394}<<<3'd2)+$signed(-{1'b0,x299})+$signed(-{2'b0,x172}<<<3'd1)+$signed({1'b0,x28})+$signed({1'b0,x221})+$signed({1'b0,x254})+$signed(-{3'b0,x207}<<<3'd2);
assign sharing22 = $signed(-{4'b0,x304}<<<3'd3)+$signed({3'b0,x305}<<<3'd2)+$signed({3'b0,x385}<<<3'd2)+$signed(-{3'b0,x49}<<<3'd2)+$signed(-{2'b0,x273}<<<3'd1)+$signed({2'b0,x418}<<<3'd1)+$signed({3'b0,x371}<<<3'd2)+$signed(-{3'b0,x35}<<<3'd2)+$signed({2'b0,x261}<<<3'd1)+$signed(-{2'b0,x85}<<<3'd1)+$signed({3'b0,x326}<<<3'd2)+$signed(-{1'b0,x86})+$signed(-{3'b0,x23}<<<3'd2)+$signed({2'b0,x199}<<<3'd1)+$signed({3'b0,x313}<<<3'd2)+$signed({3'b0,x457}<<<3'd2)+$signed(-{3'b0,x89}<<<3'd2)+$signed(-{3'b0,x41}<<<3'd2)+$signed({3'b0,x410}<<<3'd2)+$signed(-{2'b0,x249}<<<3'd1)+$signed(-{1'b0,x234})+$signed({3'b0,x155}<<<3'd2)+$signed(-{2'b0,x491}<<<3'd1)+$signed({3'b0,x300}<<<3'd2)+$signed({2'b0,x156}<<<3'd1)+$signed({3'b0,x236}<<<3'd2)+$signed({3'b0,x333}<<<3'd2)+$signed({2'b0,x269}<<<3'd1)+$signed(-{2'b0,x398}<<<3'd1)+$signed({3'b0,x287}<<<3'd2);
assign sharing23 = $signed({2'b0,x112}<<<3'd1)+$signed({2'b0,x96}<<<3'd1)+$signed({1'b0,x16})+$signed({2'b0,x352}<<<3'd1)+$signed(-{2'b0,x192}<<<3'd1)+$signed(-{1'b0,x161})+$signed(-{3'b0,x386}<<<3'd2)+$signed({2'b0,x194}<<<3'd1)+$signed({2'b0,x482}<<<3'd1)+$signed(-{3'b0,x436}<<<3'd2)+$signed({2'b0,x292}<<<3'd1)+$signed(-{3'b0,x356}<<<3'd2)+$signed({2'b0,x422}<<<3'd1)+$signed(-{1'b0,x374})+$signed({3'b0,x39}<<<3'd2)+$signed({3'b0,x375}<<<3'd2)+$signed({2'b0,x88}<<<3'd1)+$signed({2'b0,x57}<<<3'd1)+$signed({1'b0,x489})+$signed(-{2'b0,x393}<<<3'd1)+$signed({3'b0,x58}<<<3'd2)+$signed({1'b0,x442})+$signed(-{1'b0,x394})+$signed(-{3'b0,x347}<<<3'd2)+$signed({2'b0,x459}<<<3'd1)+$signed(-{1'b0,x252})+$signed(-{3'b0,x429}<<<3'd2)+$signed({3'b0,x414}<<<3'd2)+$signed(-{2'b0,x303}<<<3'd1);
assign sharing24 = $signed(-{2'b0,x128}<<<3'd1)+$signed(-{3'b0,x321}<<<3'd2)+$signed(-{3'b0,x33}<<<3'd2)+$signed({1'b0,x129})+$signed({3'b0,x290}<<<3'd2)+$signed(-{3'b0,x323}<<<3'd2)+$signed(-{2'b0,x275}<<<3'd1)+$signed(-{3'b0,x20}<<<3'd2)+$signed(-{2'b0,x388}<<<3'd1)+$signed(-{2'b0,x4}<<<3'd1)+$signed(-{3'b0,x293}<<<3'd2)+$signed(-{2'b0,x37}<<<3'd1)+$signed({2'b0,x214}<<<3'd1)+$signed({1'b0,x406})+$signed({1'b0,x6})+$signed(-{2'b0,x55}<<<3'd1)+$signed(-{1'b0,x56})+$signed(-{2'b0,x121}<<<3'd1)+$signed({1'b0,x41})+$signed(-{3'b0,x474}<<<3'd2)+$signed({2'b0,x74}<<<3'd1)+$signed(-{1'b0,x410})+$signed({2'b0,x43}<<<3'd1)+$signed(-{3'b0,x396}<<<3'd2)+$signed(-{3'b0,x124}<<<3'd2)+$signed({3'b0,x173}<<<3'd2)+$signed(-{2'b0,x109}<<<3'd1)+$signed(-{2'b0,x221}<<<3'd1)+$signed(-{1'b0,x318})+$signed({3'b0,x111}<<<3'd2);
assign sharing25 = $signed({3'b0,x224}<<<3'd2)+$signed(-{2'b0,x145}<<<3'd1)+$signed({1'b0,x193})+$signed({2'b0,x418}<<<3'd1)+$signed({2'b0,x194}<<<3'd1)+$signed(-{2'b0,x98}<<<3'd1)+$signed(-{1'b0,x19})+$signed({1'b0,x453})+$signed(-{1'b0,x245})+$signed({3'b0,x278}<<<3'd2)+$signed({3'b0,x135}<<<3'd2)+$signed({2'b0,x119}<<<3'd1)+$signed({3'b0,x344}<<<3'd2)+$signed(-{3'b0,x249}<<<3'd2)+$signed(-{1'b0,x473})+$signed(-{1'b0,x201})+$signed({3'b0,x26}<<<3'd2)+$signed({2'b0,x42}<<<3'd1)+$signed(-{1'b0,x378})+$signed({3'b0,x299}<<<3'd2)+$signed({2'b0,x395}<<<3'd1)+$signed({1'b0,x91})+$signed({3'b0,x108}<<<3'd2)+$signed({3'b0,x174}<<<3'd2)+$signed(-{2'b0,x189}<<<3'd1)+$signed({1'b0,x29})+$signed({3'b0,x158}<<<3'd2)+$signed({2'b0,x222}<<<3'd1)+$signed(-{4'b0,x463}<<<3'd3);
assign sharing26 = $signed({3'b0,x400}<<<3'd2)+$signed(-{2'b0,x272}<<<3'd1)+$signed({3'b0,x273}<<<3'd2)+$signed({2'b0,x97}<<<3'd1)+$signed({3'b0,x210}<<<3'd2)+$signed({1'b0,x2})+$signed(-{1'b0,x323})+$signed(-{1'b0,x115})+$signed(-{3'b0,x308}<<<3'd2)+$signed({3'b0,x165}<<<3'd2)+$signed({3'b0,x197}<<<3'd2)+$signed({1'b0,x229})+$signed({3'b0,x70}<<<3'd2)+$signed({3'b0,x374}<<<3'd2)+$signed({1'b0,x278})+$signed({3'b0,x40}<<<3'd2)+$signed({2'b0,x136}<<<3'd1)+$signed(-{1'b0,x472})+$signed({2'b0,x313}<<<3'd1)+$signed({3'b0,x459}<<<3'd2)+$signed(-{1'b0,x299})+$signed({3'b0,x156}<<<3'd2)+$signed(-{3'b0,x12}<<<3'd2)+$signed(-{3'b0,x461}<<<3'd2)+$signed(-{2'b0,x429}<<<3'd1)+$signed({2'b0,x222}<<<3'd1)+$signed(-{1'b0,x334})+$signed(-{2'b0,x206}<<<3'd1);
assign sharing27 = $signed(-{2'b0,x384}<<<3'd1)+$signed({1'b0,x432})+$signed({3'b0,x129}<<<3'd2)+$signed({2'b0,x257}<<<3'd1)+$signed(-{1'b0,x417})+$signed({2'b0,x50}<<<3'd1)+$signed({2'b0,x418}<<<3'd1)+$signed({2'b0,x178}<<<3'd1)+$signed(-{3'b0,x339}<<<3'd2)+$signed(-{2'b0,x99}<<<3'd1)+$signed({1'b0,x227})+$signed(-{3'b0,x483}<<<3'd2)+$signed(-{3'b0,x324}<<<3'd2)+$signed(-{2'b0,x20}<<<3'd1)+$signed({1'b0,x196})+$signed(-{3'b0,x452}<<<3'd2)+$signed(-{2'b0,x116}<<<3'd1)+$signed(-{3'b0,x38}<<<3'd2)+$signed(-{2'b0,x262}<<<3'd1)+$signed({2'b0,x231}<<<3'd1)+$signed(-{1'b0,x167})+$signed({3'b0,x57}<<<3'd2)+$signed({2'b0,x393}<<<3'd1)+$signed({2'b0,x409}<<<3'd1)+$signed(-{2'b0,x169}<<<3'd1)+$signed(-{3'b0,x426}<<<3'd2)+$signed({2'b0,x106}<<<3'd1)+$signed({1'b0,x330})+$signed(-{2'b0,x298}<<<3'd1)+$signed(-{3'b0,x428}<<<3'd2)+$signed({2'b0,x348}<<<3'd1)+$signed(-{3'b0,x349}<<<3'd2)+$signed(-{2'b0,x157}<<<3'd1)+$signed({2'b0,x495}<<<3'd1);
assign sharing28 = $signed(-{3'b0,x272}<<<3'd2)+$signed({2'b0,x96}<<<3'd1)+$signed({1'b0,x352})+$signed(-{3'b0,x0}<<<3'd2)+$signed({3'b0,x321}<<<3'd2)+$signed(-{2'b0,x160}<<<3'd1)+$signed({1'b0,x33})+$signed(-{3'b0,x481}<<<3'd2)+$signed(-{1'b0,x17})+$signed({2'b0,x434}<<<3'd1)+$signed(-{3'b0,x34}<<<3'd2)+$signed(-{1'b0,x130})+$signed(-{1'b0,x50})+$signed({3'b0,x84}<<<3'd2)+$signed({2'b0,x244}<<<3'd1)+$signed(-{3'b0,x292}<<<3'd2)+$signed(-{1'b0,x308})+$signed(-{4'b0,x181}<<<3'd3)+$signed({1'b0,x85})+$signed(-{1'b0,x165})+$signed({3'b0,x278}<<<3'd2)+$signed(-{1'b0,x230})+$signed(-{1'b0,x55})+$signed({3'b0,x328}<<<3'd2)+$signed(-{2'b0,x9}<<<3'd1)+$signed({1'b0,x265})+$signed({1'b0,x351})+$signed(-{1'b0,x25})+$signed({3'b0,x142}<<<3'd2)+$signed(-{3'b0,x396}<<<3'd2)+$signed({2'b0,x204}<<<3'd1)+$signed(-{3'b0,x220}<<<3'd2)+$signed({3'b0,x141}<<<3'd2)+$signed({3'b0,x334}<<<3'd2)+$signed({2'b0,x14}<<<3'd1)+$signed({3'b0,x399}<<<3'd2)+$signed(-{2'b0,x63}<<<3'd1)+$signed({1'b0,x15});
assign sharing29 = $signed({1'b0,x224})+$signed(-{1'b0,x304})+$signed(-{1'b0,x257})+$signed(-{1'b0,x211})+$signed(-{2'b0,x452}<<<3'd1)+$signed(-{1'b0,x180})+$signed({3'b0,x405}<<<3'd2)+$signed({2'b0,x37}<<<3'd1)+$signed({2'b0,x342}<<<3'd1)+$signed({3'b0,x119}<<<3'd2)+$signed(-{3'b0,x39}<<<3'd2)+$signed({3'b0,x248}<<<3'd2)+$signed(-{2'b0,x360}<<<3'd1)+$signed({2'b0,x122}<<<3'd1)+$signed(-{1'b0,x458})+$signed({2'b0,x459}<<<3'd1)+$signed({3'b0,x12}<<<3'd2)+$signed(-{2'b0,x332}<<<3'd1)+$signed({1'b0,x492})+$signed(-{3'b0,x253}<<<3'd2)+$signed({2'b0,x221}<<<3'd1)+$signed({3'b0,x494}<<<3'd2)+$signed({2'b0,x174}<<<3'd1)+$signed(-{3'b0,x463}<<<3'd2)+$signed({2'b0,x367}<<<3'd1);
assign sharing30 = $signed(-{1'b0,x0})+$signed({2'b0,x225}<<<3'd1)+$signed(-{1'b0,x449})+$signed(-{1'b0,x34})+$signed(-{4'b0,x37}<<<3'd3)+$signed(-{3'b0,x325}<<<3'd2)+$signed({1'b0,x232})+$signed(-{2'b0,x298}<<<3'd1)+$signed(-{1'b0,x266})+$signed(-{1'b0,x330})+$signed({3'b0,x459}<<<3'd2)+$signed(-{2'b0,x331}<<<3'd1)+$signed(-{2'b0,x107}<<<3'd1)+$signed(-{2'b0,x396}<<<3'd1)+$signed(-{2'b0,x108}<<<3'd1)+$signed(-{3'b0,x77}<<<3'd2)+$signed({1'b0,x397})+$signed({1'b0,x493})+$signed(-{3'b0,x14}<<<3'd2)+$signed({2'b0,x430}<<<3'd1)+$signed(-{1'b0,x174})+$signed(-{3'b0,x48}<<<3'd2)+$signed({3'b0,x241}<<<3'd2)+$signed(-{3'b0,x145}<<<3'd2)+$signed({1'b0,x370})+$signed({2'b0,x467}<<<3'd1)+$signed(-{1'b0,x307})+$signed(-{2'b0,x246}<<<3'd1)+$signed(-{4'b0,x55}<<<3'd3)+$signed(-{4'b0,x344}<<<3'd3)+$signed({3'b0,x280}<<<3'd2)+$signed(-{3'b0,x121}<<<3'd2)+$signed({2'b0,x25}<<<3'd1)+$signed({2'b0,x185}<<<3'd1)+$signed({1'b0,x476})+$signed(-{2'b0,x157}<<<3'd1)+$signed(-{3'b0,x127}<<<3'd2);
assign sharing31 = $signed(-{2'b0,x336}<<<3'd1)+$signed({3'b0,x273}<<<3'd2)+$signed(-{2'b0,x97}<<<3'd1)+$signed(-{2'b0,x65}<<<3'd1)+$signed({2'b0,x143}<<<3'd1)+$signed(-{2'b0,x318}<<<3'd1)+$signed({1'b0,x194})+$signed({1'b0,x434})+$signed({1'b0,x482})+$signed(-{1'b0,x146})+$signed(-{2'b0,x83}<<<3'd1)+$signed(-{3'b0,x223}<<<3'd2)+$signed({1'b0,x324})+$signed(-{2'b0,x133}<<<3'd1)+$signed(-{2'b0,x478}<<<3'd1)+$signed({2'b0,x473}<<<3'd1)+$signed({1'b0,x409})+$signed({2'b0,x474}<<<3'd1)+$signed({1'b0,x90})+$signed(-{3'b0,x11}<<<3'd2)+$signed(-{3'b0,x347}<<<3'd2)+$signed({3'b0,x332}<<<3'd2)+$signed({2'b0,x12}<<<3'd1)+$signed({2'b0,x316}<<<3'd1)+$signed({3'b0,x13}<<<3'd2)+$signed(-{3'b0,x414}<<<3'd2)+$signed({2'b0,x31}<<<3'd1)+$signed(-{3'b0,x47}<<<3'd2)+$signed({2'b0,x287}<<<3'd1)+$signed(-{1'b0,x159});
assign sharing32 = $signed(-{3'b0,x432}<<<3'd2)+$signed({2'b0,x48}<<<3'd1)+$signed({3'b0,x417}<<<3'd2)+$signed({2'b0,x241}<<<3'd1)+$signed({1'b0,x353})+$signed(-{3'b0,x177}<<<3'd2)+$signed(-{2'b0,x273}<<<3'd1)+$signed({2'b0,x130}<<<3'd1)+$signed({2'b0,x290}<<<3'd1)+$signed(-{2'b0,x18}<<<3'd1)+$signed(-{2'b0,x66}<<<3'd1)+$signed(-{1'b0,x147})+$signed(-{2'b0,x52}<<<3'd1)+$signed(-{1'b0,x164})+$signed(-{3'b0,x117}<<<3'd2)+$signed({3'b0,x326}<<<3'd2)+$signed(-{3'b0,x262}<<<3'd2)+$signed({1'b0,x134})+$signed(-{2'b0,x135}<<<3'd1)+$signed(-{2'b0,x343}<<<3'd1)+$signed(-{2'b0,x249}<<<3'd1)+$signed(-{3'b0,x138}<<<3'd2)+$signed({2'b0,x394}<<<3'd1)+$signed({3'b0,x365}<<<3'd2)+$signed(-{2'b0,x13}<<<3'd1)+$signed({1'b0,x494})+$signed({3'b0,x351}<<<3'd2)+$signed({2'b0,x223}<<<3'd1);
assign sharing33 = $signed({3'b0,x240}<<<3'd2)+$signed(-{3'b0,x384}<<<3'd2)+$signed({1'b0,x480})+$signed(-{2'b0,x80}<<<3'd1)+$signed(-{1'b0,x33})+$signed({3'b0,x50}<<<3'd2)+$signed({2'b0,x402}<<<3'd1)+$signed({1'b0,x354})+$signed(-{1'b0,x386})+$signed(-{4'b0,x99}<<<3'd3)+$signed(-{3'b0,x435}<<<3'd2)+$signed(-{3'b0,x36}<<<3'd2)+$signed({2'b0,x229}<<<3'd1)+$signed({1'b0,x197})+$signed({2'b0,x309}<<<3'd1)+$signed(-{1'b0,x5})+$signed({2'b0,x278}<<<3'd1)+$signed({2'b0,x374}<<<3'd1)+$signed({2'b0,x22}<<<3'd1)+$signed(-{1'b0,x341})+$signed(-{3'b0,x119}<<<3'd2)+$signed({1'b0,x359})+$signed(-{1'b0,x439})+$signed(-{3'b0,x383}<<<3'd2)+$signed({2'b0,x344}<<<3'd1)+$signed(-{1'b0,x424})+$signed({3'b0,x217}<<<3'd2)+$signed(-{2'b0,x345}<<<3'd1)+$signed(-{1'b0,x393})+$signed(-{2'b0,x218}<<<3'd1)+$signed(-{3'b0,x91}<<<3'd2)+$signed(-{2'b0,x491}<<<3'd1)+$signed({3'b0,x188}<<<3'd2)+$signed({2'b0,x492}<<<3'd1)+$signed(-{3'b0,x109}<<<3'd2)+$signed(-{3'b0,x382}<<<3'd2)+$signed({1'b0,x158})+$signed({3'b0,x143}<<<3'd2)+$signed(-{2'b0,x319}<<<3'd1)+$signed({1'b0,x447});
assign sharing34 = $signed({2'b0,x256}<<<3'd1)+$signed({2'b0,x320}<<<3'd1)+$signed(-{3'b0,x353}<<<3'd2)+$signed({3'b0,x66}<<<3'd2)+$signed(-{2'b0,x451}<<<3'd1)+$signed({2'b0,x388}<<<3'd1)+$signed({3'b0,x357}<<<3'd2)+$signed(-{2'b0,x423}<<<3'd1)+$signed({2'b0,x8}<<<3'd1)+$signed(-{2'b0,x264}<<<3'd1)+$signed(-{2'b0,x200}<<<3'd1)+$signed(-{1'b0,x490})+$signed(-{1'b0,x363})+$signed(-{2'b0,x12}<<<3'd1)+$signed({3'b0,x301}<<<3'd2)+$signed({3'b0,x493}<<<3'd2)+$signed(-{3'b0,x397}<<<3'd2)+$signed(-{2'b0,x237}<<<3'd1)+$signed({2'b0,x206}<<<3'd1)+$signed(-{2'b0,x334}<<<3'd1)+$signed(-{1'b0,x176})+$signed(-{3'b0,x241}<<<3'd2)+$signed(-{2'b0,x305}<<<3'd1)+$signed(-{3'b0,x114}<<<3'd2)+$signed({2'b0,x210}<<<3'd1)+$signed(-{2'b0,x178}<<<3'd1)+$signed(-{2'b0,x211}<<<3'd1)+$signed({1'b0,x147})+$signed(-{1'b0,x20})+$signed(-{2'b0,x21}<<<3'd1)+$signed(-{2'b0,x54}<<<3'd1)+$signed(-{1'b0,x342})+$signed(-{3'b0,x247}<<<3'd2)+$signed({2'b0,x343}<<<3'd1)+$signed({1'b0,x119})+$signed({3'b0,x249}<<<3'd2)+$signed({2'b0,x313}<<<3'd1)+$signed(-{3'b0,x281}<<<3'd2)+$signed(-{3'b0,x347}<<<3'd2)+$signed({3'b0,x476}<<<3'd2)+$signed({3'b0,x61}<<<3'd2)+$signed(-{3'b0,x319}<<<3'd2)+$signed({2'b0,x479}<<<3'd1);
assign sharing35 = $signed({3'b0,x384}<<<3'd2)+$signed({2'b0,x304}<<<3'd1)+$signed(-{2'b0,x81}<<<3'd1)+$signed({1'b0,x194})+$signed(-{2'b0,x275}<<<3'd1)+$signed({1'b0,x323})+$signed({2'b0,x292}<<<3'd1)+$signed({3'b0,x277}<<<3'd2)+$signed({2'b0,x405}<<<3'd1)+$signed({2'b0,x437}<<<3'd1)+$signed({1'b0,x309})+$signed(-{2'b0,x213}<<<3'd1)+$signed(-{2'b0,x182}<<<3'd1)+$signed(-{2'b0,x198}<<<3'd1)+$signed(-{2'b0,x375}<<<3'd1)+$signed(-{2'b0,x312}<<<3'd1)+$signed(-{2'b0,x377}<<<3'd1)+$signed({3'b0,x442}<<<3'd2)+$signed({2'b0,x10}<<<3'd1)+$signed({3'b0,x122}<<<3'd2)+$signed(-{3'b0,x75}<<<3'd2)+$signed(-{2'b0,x428}<<<3'd1)+$signed({3'b0,x13}<<<3'd2)+$signed({3'b0,x45}<<<3'd2)+$signed({3'b0,x205}<<<3'd2)+$signed(-{4'b0,x254}<<<3'd3)+$signed({2'b0,x303}<<<3'd1);
assign sharing36 = $signed({3'b0,x208}<<<3'd2)+$signed(-{3'b0,x113}<<<3'd2)+$signed({1'b0,x81})+$signed({1'b0,x289})+$signed(-{1'b0,x82})+$signed(-{2'b0,x387}<<<3'd1)+$signed(-{1'b0,x179})+$signed({3'b0,x84}<<<3'd2)+$signed(-{3'b0,x452}<<<3'd2)+$signed(-{1'b0,x260})+$signed(-{2'b0,x229}<<<3'd1)+$signed(-{1'b0,x357})+$signed(-{3'b0,x374}<<<3'd2)+$signed(-{3'b0,x249}<<<3'd2)+$signed({1'b0,x271})+$signed(-{2'b0,x23}<<<3'd1)+$signed({1'b0,x135})+$signed({3'b0,x88}<<<3'd2)+$signed({2'b0,x360}<<<3'd1)+$signed(-{3'b0,x488}<<<3'd2)+$signed(-{3'b0,x152}<<<3'd2)+$signed(-{4'b0,x25}<<<3'd3)+$signed({2'b0,x89}<<<3'd1)+$signed(-{2'b0,x201}<<<3'd1)+$signed(-{1'b0,x41})+$signed(-{2'b0,x105}<<<3'd1)+$signed({2'b0,x266}<<<3'd1)+$signed({2'b0,x330}<<<3'd1)+$signed(-{2'b0,x489}<<<3'd1)+$signed({3'b0,x139}<<<3'd2)+$signed({1'b0,x399})+$signed({3'b0,x379}<<<3'd2)+$signed({1'b0,x155})+$signed({2'b0,x460}<<<3'd1)+$signed({1'b0,x60})+$signed(-{2'b0,x409}<<<3'd1)+$signed({3'b0,x221}<<<3'd2)+$signed({2'b0,x413}<<<3'd1)+$signed(-{3'b0,x493}<<<3'd2)+$signed(-{3'b0,x286}<<<3'd2)+$signed({1'b0,x351});
assign sharing37 = $signed({3'b0,x464}<<<3'd2)+$signed({2'b0,x64}<<<3'd1)+$signed(-{2'b0,x48}<<<3'd1)+$signed(-{1'b0,x368})+$signed(-{1'b0,x241})+$signed(-{2'b0,x50}<<<3'd1)+$signed(-{3'b0,x340}<<<3'd2)+$signed(-{1'b0,x164})+$signed(-{2'b0,x149}<<<3'd1)+$signed(-{1'b0,x85})+$signed(-{2'b0,x102}<<<3'd1)+$signed(-{1'b0,x342})+$signed(-{3'b0,x183}<<<3'd2)+$signed(-{1'b0,x295})+$signed(-{3'b0,x120}<<<3'd2)+$signed(-{2'b0,x56}<<<3'd1)+$signed({1'b0,x168})+$signed(-{2'b0,x248}<<<3'd1)+$signed(-{2'b0,x376}<<<3'd1)+$signed({1'b0,x329})+$signed({3'b0,x186}<<<3'd2)+$signed(-{1'b0,x42})+$signed(-{1'b0,x282})+$signed(-{2'b0,x94}<<<3'd1)+$signed(-{1'b0,x491})+$signed({1'b0,x429})+$signed({2'b0,x222}<<<3'd1)+$signed({1'b0,x398})+$signed({3'b0,x367}<<<3'd2)+$signed(-{1'b0,x111});
assign sharing38 = $signed({2'b0,x416}<<<3'd1)+$signed({1'b0,x81})+$signed({1'b0,x322})+$signed({1'b0,x50})+$signed({2'b0,x195}<<<3'd1)+$signed({1'b0,x3})+$signed({2'b0,x227}<<<3'd1)+$signed({1'b0,x371})+$signed(-{1'b0,x4})+$signed({3'b0,x101}<<<3'd2)+$signed({3'b0,x22}<<<3'd2)+$signed({3'b0,x119}<<<3'd2)+$signed({2'b0,x105}<<<3'd1)+$signed({2'b0,x441}<<<3'd1)+$signed({2'b0,x249}<<<3'd1)+$signed(-{1'b0,x157})+$signed(-{2'b0,x426}<<<3'd1)+$signed({1'b0,x58})+$signed({2'b0,x459}<<<3'd1)+$signed({2'b0,x411}<<<3'd1)+$signed({3'b0,x444}<<<3'd2)+$signed(-{2'b0,x396}<<<3'd1)+$signed({1'b0,x204})+$signed({2'b0,x333}<<<3'd1)+$signed({2'b0,x365}<<<3'd1)+$signed(-{2'b0,x126}<<<3'd1);
assign sharing39 = $signed({1'b0,x256})+$signed(-{3'b0,x225}<<<3'd2)+$signed({2'b0,x321}<<<3'd1)+$signed(-{2'b0,x33}<<<3'd1)+$signed(-{1'b0,x65})+$signed({2'b0,x323}<<<3'd1)+$signed({2'b0,x261}<<<3'd1)+$signed({2'b0,x230}<<<3'd1)+$signed(-{1'b0,x38})+$signed({2'b0,x103}<<<3'd1)+$signed(-{2'b0,x39}<<<3'd1)+$signed(-{3'b0,x168}<<<3'd2)+$signed(-{3'b0,x489}<<<3'd2)+$signed(-{3'b0,x10}<<<3'd2)+$signed({2'b0,x266}<<<3'd1)+$signed(-{2'b0,x202}<<<3'd1)+$signed({3'b0,x171}<<<3'd2)+$signed(-{2'b0,x299}<<<3'd1)+$signed(-{1'b0,x75})+$signed(-{2'b0,x491}<<<3'd1)+$signed(-{1'b0,x140})+$signed(-{3'b0,x429}<<<3'd2)+$signed({2'b0,x397}<<<3'd1)+$signed(-{2'b0,x461}<<<3'd1)+$signed(-{2'b0,x398}<<<3'd1)+$signed(-{4'b0,x495}<<<3'd3)+$signed({3'b0,x175}<<<3'd2)+$signed({3'b0,x431}<<<3'd2)+$signed(-{2'b0,x239}<<<3'd1)+$signed({3'b0,x178}<<<3'd2)+$signed(-{2'b0,x434}<<<3'd1)+$signed(-{2'b0,x179}<<<3'd1)+$signed(-{1'b0,x468})+$signed(-{3'b0,x311}<<<3'd2)+$signed(-{1'b0,x23})+$signed({3'b0,x120}<<<3'd2)+$signed(-{3'b0,x376}<<<3'd2)+$signed(-{1'b0,x312})+$signed(-{1'b0,x25})+$signed(-{1'b0,x57})+$signed(-{1'b0,x313})+$signed({2'b0,x124}<<<3'd1)+$signed(-{2'b0,x61}<<<3'd1)+$signed({3'b0,x414}<<<3'd2)+$signed({1'b0,x127});
assign sharing40 = $signed(-{3'b0,x64}<<<3'd2)+$signed({2'b0,x24}<<<3'd1)+$signed({1'b0,x192})+$signed({2'b0,x152}<<<3'd1)+$signed(-{3'b0,x41}<<<3'd2)+$signed({3'b0,x42}<<<3'd2)+$signed({3'b0,x331}<<<3'd2)+$signed({2'b0,x83}<<<3'd1)+$signed(-{3'b0,x315}<<<3'd2)+$signed({4'b0,x420}<<<3'd3)+$signed(-{3'b0,x244}<<<3'd2)+$signed(-{2'b0,x396}<<<3'd1)+$signed(-{3'b0,x381}<<<3'd2)+$signed(-{2'b0,x279}<<<3'd1)+$signed(-{1'b0,x239});
assign sharing41 = $signed({1'b0,x0})+$signed(-{4'b0,x449}<<<3'd3)+$signed({3'b0,x418}<<<3'd2)+$signed({3'b0,x291}<<<3'd2)+$signed(-{3'b0,x387}<<<3'd2)+$signed(-{3'b0,x131}<<<3'd2)+$signed({3'b0,x436}<<<3'd2)+$signed(-{2'b0,x212}<<<3'd1)+$signed({2'b0,x85}<<<3'd1)+$signed(-{2'b0,x453}<<<3'd1)+$signed({4'b0,x102}<<<3'd3)+$signed(-{4'b0,x230}<<<3'd3)+$signed({2'b0,x358}<<<3'd1)+$signed(-{3'b0,x137}<<<3'd2)+$signed({2'b0,x473}<<<3'd1)+$signed(-{1'b0,x329})+$signed(-{3'b0,x410}<<<3'd2)+$signed(-{2'b0,x282}<<<3'd1)+$signed(-{1'b0,x43})+$signed({3'b0,x300}<<<3'd2)+$signed(-{3'b0,x156}<<<3'd2)+$signed(-{2'b0,x284}<<<3'd1)+$signed(-{3'b0,x29}<<<3'd2);
assign sharing42 = $signed({4'b0,x318}<<<3'd3)+$signed({1'b0,x128})+$signed({1'b0,x337})+$signed({3'b0,x18}<<<3'd2)+$signed({2'b0,x194}<<<3'd1)+$signed({3'b0,x370}<<<3'd2)+$signed(-{1'b0,x146})+$signed({2'b0,x355}<<<3'd1)+$signed(-{1'b0,x293})+$signed({2'b0,x184}<<<3'd1)+$signed({1'b0,x8})+$signed({1'b0,x377})+$signed(-{3'b0,x314}<<<3'd2)+$signed(-{1'b0,x122})+$signed(-{1'b0,x394})+$signed({3'b0,x379}<<<3'd2)+$signed({2'b0,x155}<<<3'd1)+$signed({2'b0,x315}<<<3'd1)+$signed({3'b0,x189}<<<3'd2)+$signed(-{1'b0,x13})+$signed({4'b0,x94}<<<3'd3)+$signed({3'b0,x191}<<<3'd2);
assign sharing43 = $signed({3'b0,x64}<<<3'd2)+$signed(-{3'b0,x480}<<<3'd2)+$signed(-{2'b0,x386}<<<3'd1)+$signed(-{2'b0,x242}<<<3'd1)+$signed(-{1'b0,x259})+$signed(-{1'b0,x36})+$signed(-{2'b0,x149}<<<3'd1)+$signed({3'b0,x342}<<<3'd2)+$signed(-{3'b0,x343}<<<3'd2)+$signed({2'b0,x247}<<<3'd1)+$signed(-{2'b0,x327}<<<3'd1)+$signed({1'b0,x456})+$signed(-{2'b0,x233}<<<3'd1)+$signed({1'b0,x297})+$signed({3'b0,x95}<<<3'd2)+$signed({2'b0,x271}<<<3'd1);
assign sharing44 = $signed({3'b0,x144}<<<3'd2)+$signed(-{3'b0,x160}<<<3'd2)+$signed(-{3'b0,x257}<<<3'd2)+$signed(-{1'b0,x81})+$signed(-{4'b0,x147}<<<3'd3)+$signed(-{3'b0,x244}<<<3'd2)+$signed({2'b0,x132}<<<3'd1)+$signed({2'b0,x164}<<<3'd1)+$signed(-{2'b0,x260}<<<3'd1)+$signed({3'b0,x21}<<<3'd2)+$signed({2'b0,x421}<<<3'd1)+$signed({1'b0,x5})+$signed(-{3'b0,x117}<<<3'd2)+$signed(-{1'b0,x341})+$signed({2'b0,x102}<<<3'd1)+$signed({3'b0,x313}<<<3'd2)+$signed(-{1'b0,x234})+$signed({1'b0,x141})+$signed({3'b0,x190}<<<3'd2)+$signed({2'b0,x142}<<<3'd1)+$signed({1'b0,x334});
assign sharing45 = $signed({1'b0,x240})+$signed(-{1'b0,x96})+$signed({1'b0,x49})+$signed({1'b0,x209})+$signed({1'b0,x82})+$signed(-{2'b0,x227}<<<3'd1)+$signed({2'b0,x276}<<<3'd1)+$signed({2'b0,x212}<<<3'd1)+$signed({3'b0,x69}<<<3'd2)+$signed(-{1'b0,x357})+$signed({2'b0,x470}<<<3'd1)+$signed({4'b0,x472}<<<3'd3)+$signed({2'b0,x312}<<<3'd1)+$signed({3'b0,x457}<<<3'd2)+$signed(-{2'b0,x203}<<<3'd1)+$signed(-{2'b0,x475}<<<3'd1)+$signed(-{1'b0,x267})+$signed(-{3'b0,x348}<<<3'd2)+$signed({1'b0,x444})+$signed({3'b0,x237}<<<3'd2)+$signed(-{1'b0,x303});
assign sharing46 = $signed({1'b0,x144})+$signed(-{3'b0,x433}<<<3'd2)+$signed(-{1'b0,x465})+$signed(-{3'b0,x18}<<<3'd2)+$signed(-{1'b0,x434})+$signed(-{3'b0,x324}<<<3'd2)+$signed(-{2'b0,x20}<<<3'd1)+$signed(-{1'b0,x52})+$signed(-{1'b0,x100})+$signed(-{2'b0,x325}<<<3'd1)+$signed(-{1'b0,x149})+$signed(-{4'b0,x71}<<<3'd3)+$signed(-{3'b0,x279}<<<3'd2)+$signed(-{2'b0,x471}<<<3'd1)+$signed(-{2'b0,x456}<<<3'd1)+$signed({1'b0,x185})+$signed({2'b0,x170}<<<3'd1)+$signed({2'b0,x460}<<<3'd1)+$signed(-{2'b0,x301}<<<3'd1)+$signed(-{2'b0,x317}<<<3'd1)+$signed({2'b0,x158}<<<3'd1)+$signed(-{3'b0,x495}<<<3'd2)+$signed({2'b0,x239}<<<3'd1);
assign sharing47 = $signed(-{3'b0,x400}<<<3'd2)+$signed(-{2'b0,x216}<<<3'd1)+$signed(-{3'b0,x480}<<<3'd2)+$signed({2'b0,x105}<<<3'd1)+$signed(-{2'b0,x169}<<<3'd1)+$signed(-{2'b0,x153}<<<3'd1)+$signed(-{3'b0,x146}<<<3'd2)+$signed({3'b0,x123}<<<3'd2)+$signed({3'b0,x147}<<<3'd2)+$signed({1'b0,x51})+$signed(-{2'b0,x291}<<<3'd1)+$signed(-{1'b0,x476})+$signed({3'b0,x437}<<<3'd2)+$signed(-{3'b0,x237}<<<3'd2)+$signed({1'b0,x213})+$signed(-{3'b0,x311}<<<3'd2)+$signed(-{2'b0,x310}<<<3'd1)+$signed({4'b0,x383}<<<3'd3)+$signed({3'b0,x423}<<<3'd2);
assign sharing48 = $signed(-{1'b0,x257})+$signed(-{3'b0,x146}<<<3'd2)+$signed({1'b0,x338})+$signed(-{2'b0,x291}<<<3'd1)+$signed({3'b0,x196}<<<3'd2)+$signed(-{3'b0,x255}<<<3'd2)+$signed(-{3'b0,x101}<<<3'd2)+$signed({2'b0,x287}<<<3'd1)+$signed({2'b0,x423}<<<3'd1)+$signed({3'b0,x296}<<<3'd2)+$signed({2'b0,x232}<<<3'd1)+$signed(-{3'b0,x264}<<<3'd2)+$signed(-{3'b0,x472}<<<3'd2)+$signed(-{1'b0,x408})+$signed({2'b0,x297}<<<3'd1)+$signed({3'b0,x250}<<<3'd2)+$signed({1'b0,x379})+$signed(-{2'b0,x12}<<<3'd1)+$signed({1'b0,x349})+$signed({1'b0,x190})+$signed({3'b0,x303}<<<3'd2)+$signed({2'b0,x15}<<<3'd1)+$signed(-{1'b0,x495});
assign sharing49 = $signed({3'b0,x0}<<<3'd2)+$signed({2'b0,x288}<<<3'd1)+$signed(-{3'b0,x184}<<<3'd2)+$signed(-{2'b0,x127}<<<3'd1)+$signed({1'b0,x433})+$signed({1'b0,x1})+$signed({1'b0,x57})+$signed(-{2'b0,x490}<<<3'd1)+$signed(-{2'b0,x154}<<<3'd1)+$signed(-{3'b0,x235}<<<3'd2)+$signed({1'b0,x483})+$signed(-{1'b0,x3})+$signed({2'b0,x452}<<<3'd1)+$signed(-{1'b0,x60})+$signed(-{2'b0,x165}<<<3'd1)+$signed({1'b0,x61})+$signed(-{3'b0,x270}<<<3'd2)+$signed({2'b0,x246}<<<3'd1)+$signed(-{2'b0,x295}<<<3'd1)+$signed(-{1'b0,x399});
assign sharing50 = $signed({3'b0,x16}<<<3'd2)+$signed({1'b0,x33})+$signed({3'b0,x258}<<<3'd2)+$signed(-{1'b0,x194})+$signed(-{1'b0,x18})+$signed({3'b0,x133}<<<3'd2)+$signed({2'b0,x69}<<<3'd1)+$signed({2'b0,x245}<<<3'd1)+$signed({3'b0,x438}<<<3'd2)+$signed({3'b0,x104}<<<3'd2)+$signed(-{2'b0,x473}<<<3'd1)+$signed({2'b0,x346}<<<3'd1)+$signed({1'b0,x490})+$signed(-{3'b0,x107}<<<3'd2)+$signed({2'b0,x475}<<<3'd1)+$signed({2'b0,x204}<<<3'd1)+$signed(-{1'b0,x108})+$signed({2'b0,x366}<<<3'd1)+$signed(-{1'b0,x46})+$signed(-{2'b0,x191}<<<3'd1)+$signed({1'b0,x335});
assign sharing51 = $signed(-{3'b0,x225}<<<3'd2)+$signed(-{1'b0,x305})+$signed({2'b0,x386}<<<3'd1)+$signed({2'b0,x323}<<<3'd1)+$signed({2'b0,x483}<<<3'd1)+$signed({2'b0,x436}<<<3'd1)+$signed(-{2'b0,x68}<<<3'd1)+$signed(-{2'b0,x324}<<<3'd1)+$signed({2'b0,x325}<<<3'd1)+$signed({2'b0,x182}<<<3'd1)+$signed({2'b0,x198}<<<3'd1)+$signed(-{2'b0,x294}<<<3'd1)+$signed({3'b0,x7}<<<3'd2)+$signed({2'b0,x136}<<<3'd1)+$signed({3'b0,x458}<<<3'd2)+$signed({3'b0,x251}<<<3'd2)+$signed(-{2'b0,x267}<<<3'd1)+$signed(-{3'b0,x479}<<<3'd2)+$signed({1'b0,x348})+$signed(-{1'b0,x29})+$signed(-{1'b0,x14})+$signed({3'b0,x63}<<<3'd2);
assign sharing52 = $signed(-{3'b0,x0}<<<3'd2)+$signed({2'b0,x146}<<<3'd1)+$signed({2'b0,x450}<<<3'd1)+$signed(-{2'b0,x132}<<<3'd1)+$signed({3'b0,x389}<<<3'd2)+$signed(-{2'b0,x309}<<<3'd1)+$signed(-{3'b0,x327}<<<3'd2)+$signed(-{3'b0,x295}<<<3'd2)+$signed({1'b0,x7})+$signed({1'b0,x103})+$signed(-{3'b0,x344}<<<3'd2)+$signed({1'b0,x440})+$signed({1'b0,x248})+$signed({3'b0,x282}<<<3'd2)+$signed({2'b0,x10}<<<3'd1)+$signed({1'b0,x74})+$signed(-{3'b0,x90}<<<3'd2)+$signed({1'b0,x107})+$signed(-{1'b0,x221})+$signed({3'b0,x350}<<<3'd2)+$signed({2'b0,x15}<<<3'd1);
assign sharing53 = $signed(-{3'b0,x368}<<<3'd2)+$signed({2'b0,x80}<<<3'd1)+$signed({1'b0,x176})+$signed(-{3'b0,x65}<<<3'd2)+$signed(-{3'b0,x481}<<<3'd2)+$signed({3'b0,x274}<<<3'd2)+$signed({2'b0,x3}<<<3'd1)+$signed(-{1'b0,x83})+$signed(-{3'b0,x420}<<<3'd2)+$signed(-{2'b0,x340}<<<3'd1)+$signed(-{3'b0,x37}<<<3'd2)+$signed({2'b0,x133}<<<3'd1)+$signed(-{3'b0,x118}<<<3'd2)+$signed({1'b0,x296})+$signed({3'b0,x25}<<<3'd2)+$signed({2'b0,x329}<<<3'd1)+$signed(-{3'b0,x473}<<<3'd2)+$signed(-{3'b0,x490}<<<3'd2)+$signed({3'b0,x124}<<<3'd2)+$signed({1'b0,x28})+$signed({2'b0,x173}<<<3'd1)+$signed(-{3'b0,x158}<<<3'd2)+$signed({2'b0,x286}<<<3'd1)+$signed({3'b0,x271}<<<3'd2);
assign sharing54 = $signed(-{2'b0,x304}<<<3'd1)+$signed(-{1'b0,x352})+$signed(-{3'b0,x465}<<<3'd2)+$signed({2'b0,x209}<<<3'd1)+$signed(-{2'b0,x417}<<<3'd1)+$signed(-{1'b0,x129})+$signed(-{2'b0,x450}<<<3'd1)+$signed(-{1'b0,x178})+$signed({4'b0,x371}<<<3'd3)+$signed({2'b0,x211}<<<3'd1)+$signed(-{1'b0,x131})+$signed({2'b0,x388}<<<3'd1)+$signed({2'b0,x244}<<<3'd1)+$signed(-{1'b0,x436})+$signed({2'b0,x22}<<<3'd1)+$signed(-{1'b0,x406})+$signed({2'b0,x103}<<<3'd1)+$signed(-{2'b0,x39}<<<3'd1)+$signed({2'b0,x104}<<<3'd1)+$signed(-{3'b0,x170}<<<3'd2)+$signed({2'b0,x154}<<<3'd1)+$signed({1'b0,x171})+$signed(-{1'b0,x235})+$signed(-{1'b0,x412})+$signed({1'b0,x77})+$signed({3'b0,x191}<<<3'd2)+$signed({2'b0,x479}<<<3'd1);
assign sharing55 = $signed({2'b0,x1}<<<3'd1)+$signed({1'b0,x17})+$signed(-{1'b0,x386})+$signed({2'b0,x212}<<<3'd1)+$signed({1'b0,x356})+$signed({3'b0,x293}<<<3'd2)+$signed({1'b0,x101})+$signed(-{1'b0,x438})+$signed({2'b0,x375}<<<3'd1)+$signed({2'b0,x71}<<<3'd1)+$signed(-{1'b0,x279})+$signed(-{2'b0,x440}<<<3'd1)+$signed(-{1'b0,x424})+$signed(-{3'b0,x362}<<<3'd2)+$signed({2'b0,x107}<<<3'd1)+$signed({3'b0,x444}<<<3'd2)+$signed({2'b0,x108}<<<3'd1)+$signed(-{3'b0,x76}<<<3'd2)+$signed({3'b0,x397}<<<3'd2)+$signed(-{1'b0,x301})+$signed(-{3'b0,x79}<<<3'd2)+$signed({2'b0,x175}<<<3'd1);
assign sharing56 = $signed({3'b0,x465}<<<3'd2)+$signed({2'b0,x81}<<<3'd1)+$signed(-{2'b0,x49}<<<3'd1)+$signed(-{2'b0,x404}<<<3'd1)+$signed({1'b0,x164})+$signed(-{2'b0,x36}<<<3'd1)+$signed(-{1'b0,x340})+$signed({2'b0,x453}<<<3'd1)+$signed({1'b0,x389})+$signed({2'b0,x486}<<<3'd1)+$signed(-{2'b0,x71}<<<3'd1)+$signed(-{3'b0,x312}<<<3'd2)+$signed(-{2'b0,x472}<<<3'd1)+$signed(-{3'b0,x456}<<<3'd2)+$signed({1'b0,x313})+$signed({1'b0,x329})+$signed({3'b0,x10}<<<3'd2)+$signed({2'b0,x362}<<<3'd1)+$signed({2'b0,x186}<<<3'd1)+$signed(-{3'b0,x381}<<<3'd2)+$signed(-{2'b0,x365}<<<3'd1)+$signed(-{1'b0,x317})+$signed(-{1'b0,x350});
assign sharing57 = $signed(-{1'b0,x413})+$signed({3'b0,x258}<<<3'd2)+$signed({2'b0,x163}<<<3'd1)+$signed(-{1'b0,x291})+$signed({3'b0,x388}<<<3'd2)+$signed(-{2'b0,x100}<<<3'd1)+$signed(-{1'b0,x4})+$signed(-{3'b0,x357}<<<3'd2)+$signed({1'b0,x326})+$signed({1'b0,x166})+$signed({3'b0,x183}<<<3'd2)+$signed({3'b0,x439}<<<3'd2)+$signed(-{1'b0,x102})+$signed(-{3'b0,x343}<<<3'd2)+$signed(-{3'b0,x120}<<<3'd2)+$signed(-{2'b0,x154}<<<3'd1)+$signed({1'b0,x395})+$signed({2'b0,x444}<<<3'd1)+$signed(-{1'b0,x252})+$signed({3'b0,x45}<<<3'd2)+$signed({2'b0,x205}<<<3'd1)+$signed({1'b0,x173})+$signed({2'b0,x349}<<<3'd1)+$signed(-{2'b0,x462}<<<3'd1)+$signed(-{1'b0,x110})+$signed({1'b0,x239});
assign sharing58 = $signed(-{2'b0,x448}<<<3'd1)+$signed({1'b0,x336})+$signed({2'b0,x161}<<<3'd1)+$signed({2'b0,x226}<<<3'd1)+$signed({2'b0,x354}<<<3'd1)+$signed({2'b0,x18}<<<3'd1)+$signed({4'b0,x115}<<<3'd3)+$signed({2'b0,x260}<<<3'd1)+$signed({1'b0,x244})+$signed(-{2'b0,x452}<<<3'd1)+$signed({3'b0,x133}<<<3'd2)+$signed(-{2'b0,x469}<<<3'd1)+$signed({3'b0,x7}<<<3'd2)+$signed({3'b0,x487}<<<3'd2)+$signed({3'b0,x215}<<<3'd2)+$signed({3'b0,x296}<<<3'd2)+$signed({2'b0,x280}<<<3'd1)+$signed({1'b0,x40})+$signed(-{1'b0,x344})+$signed(-{3'b0,x393}<<<3'd2)+$signed({3'b0,x218}<<<3'd2)+$signed({2'b0,x330}<<<3'd1)+$signed({3'b0,x43}<<<3'd2)+$signed({3'b0,x123}<<<3'd2)+$signed({3'b0,x364}<<<3'd2)+$signed(-{3'b0,x332}<<<3'd2)+$signed({1'b0,x156})+$signed(-{3'b0,x28}<<<3'd2)+$signed(-{1'b0,x477})+$signed(-{2'b0,x14}<<<3'd1)+$signed(-{1'b0,x286});
assign sharing59 = $signed({2'b0,x1}<<<3'd1)+$signed(-{2'b0,x49}<<<3'd1)+$signed(-{1'b0,x257})+$signed(-{2'b0,x113}<<<3'd1)+$signed({2'b0,x419}<<<3'd1)+$signed(-{1'b0,x291})+$signed(-{2'b0,x196}<<<3'd1)+$signed({2'b0,x165}<<<3'd1)+$signed(-{2'b0,x214}<<<3'd1)+$signed(-{2'b0,x151}<<<3'd1)+$signed(-{1'b0,x71})+$signed(-{2'b0,x456}<<<3'd1)+$signed({2'b0,x121}<<<3'd1)+$signed(-{2'b0,x153}<<<3'd1)+$signed({2'b0,x474}<<<3'd1)+$signed(-{1'b0,x42})+$signed({1'b0,x395})+$signed({3'b0,x93}<<<3'd2)+$signed(-{2'b0,x159}<<<3'd1)+$signed(-{1'b0,x63});
assign sharing60 = $signed({3'b0,x272}<<<3'd2)+$signed({3'b0,x304}<<<3'd2)+$signed({3'b0,x368}<<<3'd2)+$signed(-{2'b0,x488}<<<3'd1)+$signed({3'b0,x441}<<<3'd2)+$signed({2'b0,x349}<<<3'd1)+$signed(-{1'b0,x89})+$signed(-{4'b0,x318}<<<3'd3);
assign sharing61 = $signed(-{3'b0,x232}<<<3'd2)+$signed(-{2'b0,x264}<<<3'd1)+$signed({3'b0,x97}<<<3'd2)+$signed(-{2'b0,x362}<<<3'd1)+$signed(-{1'b0,x74})+$signed(-{1'b0,x186})+$signed({3'b0,x180}<<<3'd2)+$signed({2'b0,x484}<<<3'd1)+$signed({1'b0,x196})+$signed(-{3'b0,x461}<<<3'd2)+$signed({1'b0,x334})+$signed({1'b0,x422})+$signed(-{2'b0,x263}<<<3'd1);
assign sharing62 = $signed(-{3'b0,x176}<<<3'd2)+$signed({1'b0,x112})+$signed({2'b0,x258}<<<3'd1)+$signed({1'b0,x35})+$signed({2'b0,x389}<<<3'd1)+$signed({1'b0,x205})+$signed({2'b0,x381}<<<3'd1)+$signed({3'b0,x54}<<<3'd2)+$signed({2'b0,x326}<<<3'd1)+$signed(-{1'b0,x494})+$signed({3'b0,x15}<<<3'd2)+$signed({1'b0,x343});
assign sharing63 = $signed(-{1'b0,x360})+$signed(-{3'b0,x167}<<<3'd2)+$signed({1'b0,x9})+$signed({1'b0,x281})+$signed(-{3'b0,x106}<<<3'd2)+$signed({2'b0,x458}<<<3'd1)+$signed({3'b0,x163}<<<3'd2)+$signed(-{3'b0,x231}<<<3'd2)+$signed(-{2'b0,x236}<<<3'd1)+$signed(-{1'b0,x428})+$signed({2'b0,x277}<<<3'd1)+$signed(-{1'b0,x390})+$signed({1'b0,x30})+$signed({3'b0,x455}<<<3'd2);
assign sharing64 = $signed({1'b0,x240})+$signed({4'b0,x361}<<<3'd3)+$signed({3'b0,x289}<<<3'd2)+$signed(-{2'b0,x329}<<<3'd1)+$signed(-{1'b0,x233})+$signed(-{2'b0,x58}<<<3'd1)+$signed({1'b0,x346})+$signed({4'b0,x331}<<<3'd3)+$signed({3'b0,x355}<<<3'd2)+$signed({3'b0,x195}<<<3'd2)+$signed(-{3'b0,x139}<<<3'd2)+$signed(-{2'b0,x259}<<<3'd1)+$signed({3'b0,x420}<<<3'd2)+$signed(-{2'b0,x268}<<<3'd1)+$signed(-{2'b0,x188}<<<3'd1);
assign sharing65 = $signed(-{3'b0,x24}<<<3'd2)+$signed(-{2'b0,x64}<<<3'd1)+$signed({1'b0,x457})+$signed({1'b0,x449})+$signed({1'b0,x266})+$signed({2'b0,x390}<<<3'd1)+$signed(-{2'b0,x422}<<<3'd1)+$signed({2'b0,x293}<<<3'd1)+$signed(-{1'b0,x485})+$signed(-{3'b0,x94}<<<3'd2)+$signed({2'b0,x118}<<<3'd1)+$signed(-{3'b0,x327}<<<3'd2);
assign sharing66 = $signed({3'b0,x96}<<<3'd2)+$signed(-{2'b0,x144}<<<3'd1)+$signed(-{1'b0,x240})+$signed({2'b0,x361}<<<3'd1)+$signed({2'b0,x49}<<<3'd1)+$signed({2'b0,x481}<<<3'd1)+$signed({3'b0,x426}<<<3'd2)+$signed({2'b0,x313}<<<3'd1)+$signed(-{1'b0,x433})+$signed(-{3'b0,x467}<<<3'd2)+$signed({2'b0,x219}<<<3'd1)+$signed({2'b0,x300}<<<3'd1)+$signed(-{1'b0,x316})+$signed({1'b0,x269})+$signed(-{3'b0,x422}<<<3'd2)+$signed({2'b0,x238}<<<3'd1)+$signed(-{2'b0,x454}<<<3'd1);
assign sharing67 = $signed(-{3'b0,x224}<<<3'd2)+$signed({1'b0,x0})+$signed({1'b0,x264})+$signed(-{2'b0,x121}<<<3'd1)+$signed(-{2'b0,x274}<<<3'd1)+$signed({1'b0,x10})+$signed({2'b0,x52}<<<3'd1)+$signed({3'b0,x117}<<<3'd2)+$signed({2'b0,x253}<<<3'd1)+$signed(-{3'b0,x6}<<<3'd2)+$signed(-{3'b0,x278}<<<3'd2)+$signed({2'b0,x150}<<<3'd1)+$signed({2'b0,x495}<<<3'd1)+$signed({1'b0,x199});
assign sharing68 = $signed(-{2'b0,x9}<<<3'd1)+$signed({2'b0,x290}<<<3'd1)+$signed({2'b0,x466}<<<3'd1)+$signed(-{2'b0,x2}<<<3'd1)+$signed(-{1'b0,x294})+$signed({3'b0,x28}<<<3'd2)+$signed(-{2'b0,x4}<<<3'd1)+$signed(-{1'b0,x220})+$signed(-{1'b0,x44})+$signed({3'b0,x173}<<<3'd2)+$signed({2'b0,x485}<<<3'd1)+$signed(-{2'b0,x117}<<<3'd1)+$signed(-{1'b0,x61})+$signed({1'b0,x247});
assign sharing69 = $signed({2'b0,x240}<<<3'd1)+$signed(-{2'b0,x472}<<<3'd1)+$signed({2'b0,x441}<<<3'd1)+$signed({2'b0,x97}<<<3'd1)+$signed({3'b0,x354}<<<3'd2)+$signed({2'b0,x106}<<<3'd1)+$signed({2'b0,x458}<<<3'd1)+$signed(-{3'b0,x307}<<<3'd2)+$signed(-{2'b0,x243}<<<3'd1)+$signed(-{3'b0,x29}<<<3'd2)+$signed(-{3'b0,x405}<<<3'd2)+$signed(-{4'b0,x238}<<<3'd3)+$signed({3'b0,x318}<<<3'd2)+$signed({2'b0,x230}<<<3'd1)+$signed(-{3'b0,x47}<<<3'd2)+$signed(-{2'b0,x231}<<<3'd1)+$signed(-{1'b0,x143});
assign sharing70 = $signed({3'b0,x192}<<<3'd2)+$signed(-{2'b0,x368}<<<3'd1)+$signed({1'b0,x230})+$signed({2'b0,x353}<<<3'd1)+$signed({2'b0,x465}<<<3'd1)+$signed(-{2'b0,x81}<<<3'd1)+$signed(-{2'b0,x186}<<<3'd1)+$signed(-{3'b0,x187}<<<3'd2)+$signed({2'b0,x211}<<<3'd1)+$signed({2'b0,x403}<<<3'd1)+$signed({2'b0,x107}<<<3'd1)+$signed({1'b0,x62})+$signed({1'b0,x340})+$signed(-{2'b0,x117}<<<3'd1)+$signed({1'b0,x485})+$signed({1'b0,x254})+$signed(-{3'b0,x447}<<<3'd2)+$signed({2'b0,x31}<<<3'd1)+$signed(-{1'b0,x199});
assign sharing71 = $signed({2'b0,x160}<<<3'd1)+$signed(-{2'b0,x351}<<<3'd1)+$signed({2'b0,x73}<<<3'd1)+$signed(-{2'b0,x147}<<<3'd1)+$signed({2'b0,x100}<<<3'd1)+$signed(-{2'b0,x468}<<<3'd1)+$signed(-{2'b0,x134}<<<3'd1)+$signed({1'b0,x373})+$signed(-{3'b0,x22}<<<3'd2)+$signed({2'b0,x382}<<<3'd1)+$signed({2'b0,x462}<<<3'd1)+$signed({3'b0,x223}<<<3'd2)+$signed(-{2'b0,x183}<<<3'd1);
assign sharing72 = $signed({1'b0,x128})+$signed({3'b0,x153}<<<3'd2)+$signed(-{3'b0,x17}<<<3'd2)+$signed(-{2'b0,x122}<<<3'd1)+$signed({1'b0,x210})+$signed(-{2'b0,x18}<<<3'd1)+$signed({3'b0,x387}<<<3'd2)+$signed(-{3'b0,x67}<<<3'd2)+$signed({1'b0,x323})+$signed(-{2'b0,x123}<<<3'd1)+$signed({2'b0,x181}<<<3'd1)+$signed({2'b0,x341}<<<3'd1)+$signed(-{2'b0,x383}<<<3'd1);
assign sharing73 = $signed({2'b0,x384}<<<3'd1)+$signed({3'b0,x201}<<<3'd2)+$signed(-{1'b0,x257})+$signed(-{3'b0,x334}<<<3'd2)+$signed(-{3'b0,x218}<<<3'd2)+$signed({2'b0,x402}<<<3'd1)+$signed(-{2'b0,x138}<<<3'd1)+$signed({3'b0,x475}<<<3'd2)+$signed(-{3'b0,x451}<<<3'd2)+$signed({1'b0,x131})+$signed({2'b0,x452}<<<3'd1)+$signed(-{2'b0,x84}<<<3'd1)+$signed({3'b0,x421}<<<3'd2)+$signed({2'b0,x293}<<<3'd1)+$signed(-{2'b0,x197}<<<3'd1)+$signed({3'b0,x126}<<<3'd2)+$signed(-{1'b0,x278})+$signed({3'b0,x487}<<<3'd2)+$signed(-{3'b0,x222}<<<3'd2)+$signed({1'b0,x319});
assign sharing74 = $signed({3'b0,x112}<<<3'd2)+$signed({1'b0,x448})+$signed({1'b0,x238})+$signed(-{2'b0,x401}<<<3'd1)+$signed(-{3'b0,x226}<<<3'd2)+$signed({2'b0,x218}<<<3'd1)+$signed({2'b0,x139}<<<3'd1)+$signed(-{2'b0,x331}<<<3'd1)+$signed({3'b0,x100}<<<3'd2)+$signed({1'b0,x260})+$signed({3'b0,x413}<<<3'd2)+$signed({2'b0,x205}<<<3'd1)+$signed({3'b0,x477}<<<3'd2)+$signed(-{2'b0,x453}<<<3'd1)+$signed({3'b0,x494}<<<3'd2)+$signed({1'b0,x54})+$signed({2'b0,x391}<<<3'd1)+$signed(-{1'b0,x479});
assign sharing75 = $signed({1'b0,x160})+$signed({3'b0,x369}<<<3'd2)+$signed({2'b0,x281}<<<3'd1)+$signed(-{1'b0,x161})+$signed(-{1'b0,x113})+$signed({2'b0,x410}<<<3'd1)+$signed(-{1'b0,x474})+$signed({3'b0,x395}<<<3'd2)+$signed({3'b0,x147}<<<3'd2)+$signed(-{3'b0,x363}<<<3'd2)+$signed(-{2'b0,x291}<<<3'd1)+$signed({3'b0,x108}<<<3'd2)+$signed(-{2'b0,x69}<<<3'd1)+$signed({3'b0,x383}<<<3'd2)+$signed({2'b0,x487}<<<3'd1)+$signed({1'b0,x351});
assign sharing76 = $signed(-{3'b0,x144}<<<3'd2)+$signed({2'b0,x32}<<<3'd1)+$signed(-{2'b0,x328}<<<3'd1)+$signed({1'b0,x97})+$signed(-{3'b0,x434}<<<3'd2)+$signed(-{3'b0,x226}<<<3'd2)+$signed(-{2'b0,x485}<<<3'd1)+$signed(-{2'b0,x125}<<<3'd1)+$signed({1'b0,x350})+$signed(-{2'b0,x415}<<<3'd1)+$signed({1'b0,x191});
assign sharing77 = $signed(-{2'b0,x224}<<<3'd1)+$signed(-{4'b0,x129}<<<3'd3)+$signed({1'b0,x49})+$signed(-{3'b0,x258}<<<3'd2)+$signed(-{1'b0,x274})+$signed({3'b0,x100}<<<3'd2)+$signed({2'b0,x356}<<<3'd1)+$signed({1'b0,x324})+$signed({2'b0,x308}<<<3'd1)+$signed(-{2'b0,x404}<<<3'd1)+$signed(-{1'b0,x276})+$signed(-{1'b0,x471})+$signed(-{3'b0,x168}<<<3'd2)+$signed(-{2'b0,x440}<<<3'd1)+$signed(-{3'b0,x233}<<<3'd2)+$signed(-{2'b0,x425}<<<3'd1)+$signed(-{3'b0,x26}<<<3'd2)+$signed(-{3'b0,x203}<<<3'd2)+$signed({1'b0,x187})+$signed({1'b0,x267})+$signed({3'b0,x140}<<<3'd2)+$signed(-{1'b0,x123})+$signed(-{2'b0,x44}<<<3'd1)+$signed(-{1'b0,x95});
assign sharing78 = $signed({2'b0,x464}<<<3'd1)+$signed(-{2'b0,x177}<<<3'd1)+$signed(-{3'b0,x242}<<<3'd2)+$signed(-{2'b0,x146}<<<3'd1)+$signed({1'b0,x127})+$signed({2'b0,x52}<<<3'd1)+$signed({2'b0,x436}<<<3'd1)+$signed(-{4'b0,x469}<<<3'd3)+$signed(-{1'b0,x479})+$signed(-{2'b0,x374}<<<3'd1)+$signed(-{1'b0,x310})+$signed({3'b0,x23}<<<3'd2)+$signed(-{3'b0,x72}<<<3'd2)+$signed(-{3'b0,x330}<<<3'd2)+$signed({1'b0,x58})+$signed({3'b0,x316}<<<3'd2)+$signed({2'b0,x412}<<<3'd1)+$signed(-{2'b0,x397}<<<3'd1)+$signed({1'b0,x157})+$signed(-{3'b0,x430}<<<3'd2)+$signed(-{3'b0,x383}<<<3'd2)+$signed({1'b0,x31});
assign sharing79 = $signed({2'b0,x256}<<<3'd1)+$signed({1'b0,x336})+$signed(-{3'b0,x409}<<<3'd2)+$signed({3'b0,x482}<<<3'd2)+$signed({2'b0,x450}<<<3'd1)+$signed({2'b0,x370}<<<3'd1)+$signed({4'b0,x435}<<<3'd3)+$signed(-{2'b0,x315}<<<3'd1)+$signed({1'b0,x284})+$signed({3'b0,x261}<<<3'd2)+$signed(-{2'b0,x38}<<<3'd1)+$signed({3'b0,x143}<<<3'd2)+$signed({2'b0,x487}<<<3'd1);
assign sharing80 = $signed(-{1'b0,x368})+$signed({2'b0,x337}<<<3'd1)+$signed({3'b0,x186}<<<3'd2)+$signed({1'b0,x106})+$signed({3'b0,x43}<<<3'd2)+$signed({2'b0,x227}<<<3'd1)+$signed(-{2'b0,x19}<<<3'd1)+$signed(-{3'b0,x261}<<<3'd2)+$signed(-{1'b0,x310})+$signed({3'b0,x407}<<<3'd2);
assign sharing81 = $signed(-{3'b0,x280}<<<3'd2)+$signed(-{2'b0,x428}<<<3'd1)+$signed(-{2'b0,x252}<<<3'd1)+$signed({2'b0,x329}<<<3'd1)+$signed(-{1'b0,x31})+$signed({1'b0,x35});
assign sharing82 = $signed({3'b0,x240}<<<3'd2)+$signed({2'b0,x32}<<<3'd1)+$signed(-{3'b0,x353}<<<3'd2)+$signed(-{1'b0,x209})+$signed(-{2'b0,x399}<<<3'd1)+$signed(-{2'b0,x237}<<<3'd1)+$signed({2'b0,x342}<<<3'd1)+$signed(-{2'b0,x351}<<<3'd1);
assign sharing83 = $signed(-{1'b0,x408})+$signed({2'b0,x170}<<<3'd1)+$signed(-{2'b0,x282}<<<3'd1)+$signed(-{1'b0,x450})+$signed(-{3'b0,x331}<<<3'd2)+$signed(-{1'b0,x340})+$signed({3'b0,x222}<<<3'd2)+$signed(-{1'b0,x206})+$signed(-{2'b0,x183}<<<3'd1);
assign sharing84 = $signed(-{4'b0,x280}<<<3'd3)+$signed({2'b0,x240}<<<3'd1)+$signed(-{1'b0,x120})+$signed(-{4'b0,x217}<<<3'd3)+$signed({1'b0,x482})+$signed({3'b0,x44}<<<3'd2)+$signed({3'b0,x277}<<<3'd2)+$signed(-{2'b0,x30}<<<3'd1)+$signed({2'b0,x71}<<<3'd1)+$signed(-{1'b0,x175});
assign sharing85 = $signed(-{3'b0,x320}<<<3'd2)+$signed(-{3'b0,x105}<<<3'd2)+$signed(-{2'b0,x361}<<<3'd1)+$signed(-{3'b0,x164}<<<3'd2)+$signed({2'b0,x77}<<<3'd1)+$signed(-{2'b0,x45}<<<3'd1)+$signed(-{3'b0,x182}<<<3'd2)+$signed(-{1'b0,x398})+$signed(-{4'b0,x311}<<<3'd3);
assign sharing86 = $signed({2'b0,x6}<<<3'd1)+$signed(-{1'b0,x89})+$signed({3'b0,x490}<<<3'd2)+$signed(-{3'b0,x234}<<<3'd2)+$signed(-{3'b0,x435}<<<3'd2)+$signed({2'b0,x427}<<<3'd1)+$signed({3'b0,x196}<<<3'd2)+$signed(-{2'b0,x20}<<<3'd1)+$signed({1'b0,x76})+$signed(-{2'b0,x92}<<<3'd1)+$signed({2'b0,x245}<<<3'd1)+$signed({1'b0,x213})+$signed({2'b0,x150}<<<3'd1)+$signed({1'b0,x214});
assign sharing87 = $signed({3'b0,x292}<<<3'd2)+$signed(-{2'b0,x300}<<<3'd1)+$signed(-{2'b0,x364}<<<3'd1)+$signed(-{1'b0,x21})+$signed({4'b0,x455}<<<3'd3)+$signed(-{1'b0,x243});
assign sharing88 = $signed({4'b0,x408}<<<3'd3)+$signed(-{3'b0,x305}<<<3'd2)+$signed(-{2'b0,x490}<<<3'd1)+$signed(-{3'b0,x27}<<<3'd2)+$signed(-{1'b0,x469})+$signed({3'b0,x69}<<<3'd2)+$signed({2'b0,x333}<<<3'd1)+$signed({1'b0,x53})+$signed(-{3'b0,x285}<<<3'd2)+$signed(-{1'b0,x134});
assign sharing89 = $signed({2'b0,x112}<<<3'd1)+$signed(-{2'b0,x72}<<<3'd1)+$signed({2'b0,x385}<<<3'd1)+$signed(-{2'b0,x482}<<<3'd1)+$signed({4'b0,x115}<<<3'd3)+$signed(-{3'b0,x223}<<<3'd2)+$signed({2'b0,x187}<<<3'd1)+$signed({3'b0,x389}<<<3'd2)+$signed({3'b0,x206}<<<3'd2)+$signed({3'b0,x335}<<<3'd2);
assign sharing90 = $signed(-{3'b0,x129}<<<3'd2)+$signed({1'b0,x321})+$signed({2'b0,x394}<<<3'd1)+$signed({2'b0,x338}<<<3'd1)+$signed(-{1'b0,x114})+$signed({3'b0,x403}<<<3'd2)+$signed(-{4'b0,x388}<<<3'd3)+$signed(-{3'b0,x100}<<<3'd2)+$signed({3'b0,x53}<<<3'd2)+$signed(-{3'b0,x109}<<<3'd2)+$signed({3'b0,x255}<<<3'd2)+$signed(-{1'b0,x463});
assign sharing91 = $signed(-{1'b0,x448})+$signed(-{2'b0,x17}<<<3'd1)+$signed({3'b0,x290}<<<3'd2)+$signed({2'b0,x250}<<<3'd1)+$signed({2'b0,x442}<<<3'd1)+$signed(-{3'b0,x308}<<<3'd2)+$signed({3'b0,x86}<<<3'd2)+$signed(-{3'b0,x262}<<<3'd2);
assign sharing92 = $signed(-{2'b0,x200}<<<3'd1)+$signed({3'b0,x425}<<<3'd2)+$signed({2'b0,x433}<<<3'd1)+$signed(-{3'b0,x366}<<<3'd2)+$signed(-{2'b0,x188}<<<3'd1)+$signed(-{2'b0,x140}<<<3'd1)+$signed(-{2'b0,x164}<<<3'd1)+$signed(-{3'b0,x5}<<<3'd2)+$signed({1'b0,x253})+$signed(-{3'b0,x46}<<<3'd2)+$signed(-{1'b0,x246})+$signed(-{2'b0,x463}<<<3'd1);
assign sharing93 = $signed(-{1'b0,x109})+$signed({3'b0,x345}<<<3'd2)+$signed({2'b0,x217}<<<3'd1)+$signed({3'b0,x33}<<<3'd2)+$signed({2'b0,x277}<<<3'd1)+$signed(-{1'b0,x405})+$signed(-{2'b0,x101}<<<3'd1)+$signed(-{1'b0,x170})+$signed({2'b0,x251}<<<3'd1);
assign sharing94 = $signed(-{1'b0,x440})+$signed(-{1'b0,x322})+$signed(-{3'b0,x443}<<<3'd2)+$signed(-{3'b0,x324}<<<3'd2)+$signed({4'b0,x277}<<<3'd3)+$signed({1'b0,x77})+$signed({4'b0,x478}<<<3'd3)+$signed({3'b0,x462}<<<3'd2)+$signed({2'b0,x390}<<<3'd1)+$signed({3'b0,x246}<<<3'd2)+$signed({3'b0,x191}<<<3'd2);
assign sharing95 = $signed(-{4'b0,x377}<<<3'd3)+$signed(-{3'b0,x179}<<<3'd2)+$signed(-{2'b0,x459}<<<3'd1)+$signed(-{1'b0,x46})+$signed(-{2'b0,x172}<<<3'd1)+$signed({1'b0,x100})+$signed({4'b0,x485}<<<3'd3)+$signed(-{2'b0,x292}<<<3'd1)+$signed({2'b0,x149}<<<3'd1)+$signed(-{1'b0,x477})+$signed({1'b0,x94})+$signed(-{3'b0,x495}<<<3'd2);
assign sharing96 = $signed(-{2'b0,x104}<<<3'd1)+$signed(-{2'b0,x262}<<<3'd1)+$signed({3'b0,x97}<<<3'd2)+$signed(-{3'b0,x299}<<<3'd2)+$signed(-{1'b0,x83})+$signed(-{1'b0,x175})+$signed({2'b0,x22}<<<3'd1)+$signed({1'b0,x135});
assign sharing97 = $signed({3'b0,x288}<<<3'd2)+$signed({3'b0,x416}<<<3'd2)+$signed({1'b0,x441})+$signed({3'b0,x394}<<<3'd2)+$signed(-{3'b0,x322}<<<3'd2)+$signed(-{3'b0,x386}<<<3'd2)+$signed({4'b0,x403}<<<3'd3)+$signed(-{2'b0,x3}<<<3'd1)+$signed({3'b0,x92}<<<3'd2)+$signed({2'b0,x348}<<<3'd1)+$signed({1'b0,x132})+$signed(-{1'b0,x300})+$signed(-{3'b0,x341}<<<3'd2)+$signed(-{1'b0,x414})+$signed({3'b0,x359}<<<3'd2);
assign sharing98 = $signed(-{2'b0,x288}<<<3'd1)+$signed(-{4'b0,x17}<<<3'd3)+$signed(-{4'b0,x338}<<<3'd3)+$signed({3'b0,x115}<<<3'd2)+$signed(-{3'b0,x435}<<<3'd2)+$signed(-{4'b0,x53}<<<3'd3)+$signed({3'b0,x181}<<<3'd2)+$signed(-{3'b0,x262}<<<3'd2)+$signed({1'b0,x6})+$signed({2'b0,x74}<<<3'd1)+$signed(-{3'b0,x59}<<<3'd2)+$signed(-{3'b0,x316}<<<3'd2)+$signed(-{1'b0,x332})+$signed({4'b0,x253}<<<3'd3)+$signed(-{3'b0,x77}<<<3'd2)+$signed(-{3'b0,x30}<<<3'd2)+$signed({2'b0,x207}<<<3'd1);
assign sharing99 = $signed({4'b0,x104}<<<3'd3)+$signed(-{3'b0,x360}<<<3'd2)+$signed(-{1'b0,x232})+$signed(-{3'b0,x217}<<<3'd2)+$signed({1'b0,x481})+$signed(-{3'b0,x395}<<<3'd2)+$signed(-{3'b0,x412}<<<3'd2)+$signed({3'b0,x469}<<<3'd2)+$signed({3'b0,x165}<<<3'd2)+$signed({2'b0,x190}<<<3'd1)+$signed(-{2'b0,x391}<<<3'd1);
assign sharing100 = $signed({2'b0,x392}<<<3'd1)+$signed(-{2'b0,x425}<<<3'd1)+$signed({3'b0,x443}<<<3'd2)+$signed({3'b0,x51}<<<3'd2)+$signed({2'b0,x83}<<<3'd1)+$signed(-{1'b0,x451});
assign sharing101 = $signed(-{3'b0,x160}<<<3'd2)+$signed({2'b0,x148}<<<3'd1)+$signed(-{1'b0,x272})+$signed(-{2'b0,x13}<<<3'd1)+$signed(-{4'b0,x118}<<<3'd3)+$signed({3'b0,x74}<<<3'd2)+$signed(-{1'b0,x246});
assign sharing102 = $signed({2'b0,x319}<<<3'd1)+$signed({3'b0,x169}<<<3'd2)+$signed({1'b0,x133})+$signed({1'b0,x341})+$signed({3'b0,x390}<<<3'd2)+$signed({2'b0,x347}<<<3'd1)+$signed({1'b0,x423});
assign sharing103 = $signed({2'b0,x56}<<<3'd1)+$signed(-{1'b0,x288})+$signed(-{3'b0,x98}<<<3'd2)+$signed({2'b0,x99}<<<3'd1)+$signed(-{3'b0,x116}<<<3'd2)+$signed(-{1'b0,x324})+$signed({2'b0,x37}<<<3'd1)+$signed({1'b0,x165});
assign sharing104 = $signed(-{4'b0,x416}<<<3'd3)+$signed({1'b0,x136})+$signed(-{1'b0,x360})+$signed(-{1'b0,x178})+$signed({1'b0,x245})+$signed(-{3'b0,x358}<<<3'd2)+$signed({2'b0,x62}<<<3'd1)+$signed({1'b0,x462})+$signed(-{2'b0,x367}<<<3'd1);
assign sharing105 = $signed(-{3'b0,x348}<<<3'd2)+$signed({1'b0,x20})+$signed({4'b0,x189}<<<3'd3)+$signed(-{1'b0,x401})+$signed({2'b0,x426}<<<3'd1)+$signed(-{1'b0,x306})+$signed({3'b0,x219}<<<3'd2);
assign sharing106 = $signed(-{1'b0,x466})+$signed({1'b0,x48})+$signed(-{3'b0,x431}<<<3'd2)+$signed({2'b0,x11}<<<3'd1);
assign sharing107 = $signed(-{2'b0,x120}<<<3'd1)+$signed(-{3'b0,x449}<<<3'd2)+$signed(-{1'b0,x226})+$signed(-{2'b0,x131}<<<3'd1)+$signed(-{2'b0,x451}<<<3'd1)+$signed(-{1'b0,x460})+$signed(-{4'b0,x93}<<<3'd3)+$signed(-{3'b0,x197}<<<3'd2)+$signed(-{2'b0,x301}<<<3'd1)+$signed({2'b0,x350}<<<3'd1)+$signed({1'b0,x118})+$signed({3'b0,x295}<<<3'd2);
assign sharing108 = $signed({3'b0,x464}<<<3'd2)+$signed({1'b0,x152})+$signed({1'b0,x212})+$signed({1'b0,x172})+$signed({1'b0,x348})+$signed(-{2'b0,x69}<<<3'd1)+$signed(-{3'b0,x274}<<<3'd2)+$signed(-{2'b0,x155}<<<3'd1)+$signed({1'b0,x491});
assign sharing109 = $signed({2'b0,x377}<<<3'd1)+$signed({2'b0,x306}<<<3'd1)+$signed(-{3'b0,x374}<<<3'd2)+$signed({2'b0,x139}<<<3'd1)+$signed(-{3'b0,x484}<<<3'd2)+$signed(-{2'b0,x5}<<<3'd1)+$signed(-{3'b0,x142}<<<3'd2)+$signed(-{2'b0,x191}<<<3'd1);
assign sharing110 = $signed({1'b0,x32})+$signed(-{1'b0,x185})+$signed({2'b0,x74}<<<3'd1)+$signed({2'b0,x419}<<<3'd1)+$signed({2'b0,x35}<<<3'd1)+$signed(-{2'b0,x203}<<<3'd1)+$signed({2'b0,x172}<<<3'd1)+$signed({2'b0,x412}<<<3'd1)+$signed({1'b0,x124})+$signed(-{1'b0,x492})+$signed(-{2'b0,x407}<<<3'd1);
assign sharing111 = $signed({3'b0,x288}<<<3'd2)+$signed(-{3'b0,x372}<<<3'd2)+$signed(-{1'b0,x444})+$signed(-{3'b0,x306}<<<3'd2)+$signed(-{2'b0,x158}<<<3'd1)+$signed(-{3'b0,x319}<<<3'd2);
assign sharing112 = $signed(-{2'b0,x168}<<<3'd1)+$signed(-{1'b0,x321})+$signed({2'b0,x362}<<<3'd1)+$signed({1'b0,x98})+$signed({3'b0,x179}<<<3'd2)+$signed({3'b0,x411}<<<3'd2)+$signed(-{2'b0,x243}<<<3'd1)+$signed({4'b0,x444}<<<3'd3)+$signed(-{2'b0,x252}<<<3'd1)+$signed({3'b0,x365}<<<3'd2)+$signed(-{3'b0,x261}<<<3'd2)+$signed({1'b0,x333})+$signed({2'b0,x455}<<<3'd1);
assign sharing113 = $signed({1'b0,x39})+$signed({2'b0,x60}<<<3'd1)+$signed({1'b0,x242})+$signed({1'b0,x318});
assign sharing114 = $signed(-{3'b0,x80}<<<3'd2)+$signed(-{3'b0,x200}<<<3'd2)+$signed(-{3'b0,x264}<<<3'd2)+$signed(-{1'b0,x412})+$signed(-{3'b0,x207}<<<3'd2)+$signed({2'b0,x271}<<<3'd1);
assign sharing115 = $signed({3'b0,x16}<<<3'd2)+$signed(-{1'b0,x425})+$signed({3'b0,x2}<<<3'd2)+$signed({2'b0,x42}<<<3'd1)+$signed({3'b0,x155}<<<3'd2)+$signed(-{1'b0,x283})+$signed(-{4'b0,x356}<<<3'd3)+$signed({3'b0,x38}<<<3'd2)+$signed({2'b0,x294}<<<3'd1)+$signed(-{1'b0,x486})+$signed(-{3'b0,x103}<<<3'd2);
assign sharing116 = $signed(-{3'b0,x56}<<<3'd2)+$signed({4'b0,x370}<<<3'd3)+$signed(-{4'b0,x122}<<<3'd3)+$signed({2'b0,x250}<<<3'd1)+$signed({1'b0,x26})+$signed({2'b0,x339}<<<3'd1)+$signed({1'b0,x124})+$signed(-{4'b0,x293}<<<3'd3)+$signed(-{1'b0,x182})+$signed(-{1'b0,x79});
assign sharing117 = $signed({2'b0,x408}<<<3'd1)+$signed({4'b0,x25}<<<3'd3)+$signed({2'b0,x257}<<<3'd1)+$signed({1'b0,x361})+$signed({3'b0,x10}<<<3'd2)+$signed(-{1'b0,x154})+$signed({3'b0,x411}<<<3'd2)+$signed({2'b0,x126}<<<3'd1)+$signed({3'b0,x463}<<<3'd2);
assign sharing118 = $signed({1'b0,x280})+$signed({2'b0,x433}<<<3'd1)+$signed(-{2'b0,x457}<<<3'd1)+$signed(-{1'b0,x246})+$signed({1'b0,x188})+$signed({3'b0,x333}<<<3'd2)+$signed({2'b0,x373}<<<3'd1)+$signed(-{1'b0,x270})+$signed({2'b0,x87}<<<3'd1)+$signed(-{1'b0,x335});
assign sharing119 = $signed({3'b0,x344}<<<3'd2)+$signed({3'b0,x112}<<<3'd2)+$signed({3'b0,x417}<<<3'd2)+$signed({2'b0,x489}<<<3'd1)+$signed({1'b0,x273})+$signed({3'b0,x474}<<<3'd2)+$signed({1'b0,x354})+$signed({3'b0,x99}<<<3'd2)+$signed({1'b0,x11})+$signed({3'b0,x172}<<<3'd2)+$signed({1'b0,x372})+$signed({4'b0,x117}<<<3'd3)+$signed({3'b0,x390}<<<3'd2)+$signed({2'b0,x382}<<<3'd1)+$signed(-{4'b0,x111}<<<3'd3);
assign sharing120 = $signed(-{3'b0,x257}<<<3'd2)+$signed(-{2'b0,x449}<<<3'd1)+$signed(-{1'b0,x437})+$signed({1'b0,x68})+$signed({2'b0,x125}<<<3'd1)+$signed(-{2'b0,x93}<<<3'd1)+$signed(-{3'b0,x454}<<<3'd2)+$signed(-{1'b0,x159});
assign sharing121 = $signed(-{1'b0,x202})+$signed({1'b0,x40})+$signed({3'b0,x445}<<<3'd2)+$signed({2'b0,x334}<<<3'd1)+$signed(-{1'b0,x70})+$signed({1'b0,x459});
assign sharing122 = $signed({2'b0,x456}<<<3'd1)+$signed(-{2'b0,x128}<<<3'd1)+$signed(-{1'b0,x59})+$signed(-{3'b0,x377}<<<3'd2)+$signed(-{2'b0,x163}<<<3'd1)+$signed({1'b0,x347});
assign sharing123 = $signed({3'b0,x404}<<<3'd2)+$signed({1'b0,x320})+$signed(-{3'b0,x117}<<<3'd2)+$signed(-{1'b0,x473})+$signed(-{3'b0,x194}<<<3'd2)+$signed(-{1'b0,x78});
assign sharing124 = $signed(-{2'b0,x164}<<<3'd1)+$signed({1'b0,x384})+$signed(-{4'b0,x97}<<<3'd3)+$signed({2'b0,x413}<<<3'd1)+$signed({3'b0,x102}<<<3'd2)+$signed(-{1'b0,x262});
assign sharing125 = $signed({4'b0,x480}<<<3'd3)+$signed({3'b0,x407}<<<3'd2)+$signed(-{3'b0,x297}<<<3'd2)+$signed({2'b0,x137}<<<3'd1)+$signed({2'b0,x162}<<<3'd1)+$signed(-{2'b0,x67}<<<3'd1)+$signed({4'b0,x236}<<<3'd3)+$signed(-{3'b0,x84}<<<3'd2)+$signed({2'b0,x116}<<<3'd1)+$signed(-{3'b0,x36}<<<3'd2)+$signed(-{2'b0,x101}<<<3'd1)+$signed({3'b0,x391}<<<3'd2);
assign sharing126 = $signed({3'b0,x64}<<<3'd2)+$signed({2'b0,x224}<<<3'd1)+$signed({3'b0,x209}<<<3'd2)+$signed({2'b0,x145}<<<3'd1)+$signed({1'b0,x121})+$signed({3'b0,x227}<<<3'd2)+$signed(-{1'b0,x251})+$signed({3'b0,x108}<<<3'd2)+$signed(-{2'b0,x189}<<<3'd1)+$signed(-{2'b0,x94}<<<3'd1)+$signed(-{1'b0,x223});
assign sharing127 = $signed({3'b0,x378}<<<3'd2)+$signed(-{2'b0,x264}<<<3'd1)+$signed(-{1'b0,x276});
assign sharing128 = $signed({2'b0,x321}<<<3'd1)+$signed({2'b0,x445}<<<3'd1)+$signed({3'b0,x458}<<<3'd2)+$signed({1'b0,x42})+$signed({3'b0,x471}<<<3'd2);
assign sharing129 = $signed({2'b0,x144}<<<3'd1)+$signed({1'b0,x44})+$signed({1'b0,x52})+$signed(-{1'b0,x224})+$signed(-{1'b0,x261})+$signed(-{3'b0,x466}<<<3'd2)+$signed({3'b0,x410}<<<3'd2)+$signed(-{2'b0,x267}<<<3'd1)+$signed({2'b0,x303}<<<3'd1);
assign sharing130 = $signed({4'b0,x400}<<<3'd3)+$signed(-{2'b0,x432}<<<3'd1)+$signed({1'b0,x177})+$signed(-{1'b0,x189})+$signed({3'b0,x166}<<<3'd2)+$signed(-{2'b0,x374}<<<3'd1)+$signed(-{1'b0,x370})+$signed({3'b0,x15}<<<3'd2)+$signed({1'b0,x399});
assign sharing131 = $signed({1'b0,x480})+$signed(-{2'b0,x185}<<<3'd1)+$signed(-{1'b0,x145})+$signed(-{2'b0,x90}<<<3'd1)+$signed(-{3'b0,x383}<<<3'd2)+$signed({2'b0,x223}<<<3'd1);
assign sharing132 = $signed(-{2'b0,x215}<<<3'd1)+$signed(-{2'b0,x239}<<<3'd1)+$signed({3'b0,x385}<<<3'd2)+$signed({3'b0,x329}<<<3'd2)+$signed({1'b0,x481})+$signed({3'b0,x181}<<<3'd2)+$signed({3'b0,x437}<<<3'd2)+$signed(-{1'b0,x177})+$signed({2'b0,x99}<<<3'd1);
assign sharing133 = $signed({4'b0,x365}<<<3'd3)+$signed(-{1'b0,x113})+$signed(-{1'b0,x150})+$signed({1'b0,x138})+$signed({3'b0,x335}<<<3'd2)+$signed({2'b0,x411}<<<3'd1);
assign sharing134 = $signed({3'b0,x128}<<<3'd2)+$signed(-{3'b0,x456}<<<3'd2)+$signed(-{1'b0,x200})+$signed({3'b0,x49}<<<3'd2)+$signed({1'b0,x266})+$signed({3'b0,x19}<<<3'd2)+$signed({2'b0,x51}<<<3'd1)+$signed({1'b0,x211})+$signed(-{1'b0,x283})+$signed(-{2'b0,x406}<<<3'd1)+$signed(-{3'b0,x63}<<<3'd2);
assign sharing135 = $signed(-{3'b0,x190}<<<3'd2)+$signed(-{2'b0,x430}<<<3'd1)+$signed(-{3'b0,x11}<<<3'd2)+$signed(-{2'b0,x86}<<<3'd1);
assign sharing136 = $signed(-{4'b0,x284}<<<3'd3)+$signed(-{2'b0,x494}<<<3'd1)+$signed({2'b0,x152}<<<3'd1)+$signed({3'b0,x205}<<<3'd2)+$signed(-{2'b0,x465}<<<3'd1)+$signed({3'b0,x238}<<<3'd2)+$signed({2'b0,x302}<<<3'd1)+$signed({2'b0,x435}<<<3'd1)+$signed(-{2'b0,x279}<<<3'd1);
assign sharing137 = $signed(-{1'b0,x56})+$signed(-{4'b0,x113}<<<3'd3)+$signed({3'b0,x339}<<<3'd2)+$signed(-{3'b0,x203}<<<3'd2)+$signed({3'b0,x12}<<<3'd2)+$signed(-{3'b0,x260}<<<3'd2)+$signed(-{3'b0,x213}<<<3'd2)+$signed(-{1'b0,x47});
assign sharing138 = $signed(-{2'b0,x486}<<<3'd1)+$signed({3'b0,x355}<<<3'd2)+$signed({2'b0,x299}<<<3'd1);
assign sharing139 = $signed(-{3'b0,x468}<<<3'd2)+$signed(-{2'b0,x122}<<<3'd1)+$signed({1'b0,x92})+$signed({1'b0,x281})+$signed(-{2'b0,x410}<<<3'd1);
assign sharing140 = $signed({3'b0,x114}<<<3'd2)+$signed(-{1'b0,x418})+$signed({1'b0,x155})+$signed({2'b0,x147}<<<3'd1)+$signed({1'b0,x271});
assign sharing141 = $signed({2'b0,x198}<<<3'd1)+$signed({3'b0,x307}<<<3'd2)+$signed({3'b0,x301}<<<3'd2);
assign sharing142 = $signed(-{1'b0,x328})+$signed({2'b0,x173}<<<3'd1)+$signed({1'b0,x413})+$signed(-{2'b0,x429}<<<3'd1)+$signed(-{1'b0,x458})+$signed(-{1'b0,x431});
assign sharing143 = $signed(-{2'b0,x48}<<<3'd1)+$signed(-{1'b0,x398})+$signed({1'b0,x315});
assign sharing144 = $signed({3'b0,x76}<<<3'd2)+$signed({3'b0,x25}<<<3'd2)+$signed({4'b0,x362}<<<3'd3)+$signed(-{3'b0,x422}<<<3'd2)+$signed({3'b0,x367}<<<3'd2);
assign sharing145 = $signed({3'b0,x169}<<<3'd2)+$signed(-{3'b0,x229}<<<3'd2)+$signed({1'b0,x345})+$signed({3'b0,x86}<<<3'd2)+$signed({1'b0,x34});
assign sharing146 = $signed({1'b0,x256})+$signed({4'b0,x273}<<<3'd3)+$signed(-{2'b0,x345}<<<3'd1)+$signed(-{3'b0,x246}<<<3'd2)+$signed({4'b0,x375}<<<3'd3)+$signed(-{1'b0,x443});
assign sharing147 = $signed({3'b0,x432}<<<3'd2)+$signed(-{2'b0,x344}<<<3'd1)+$signed({4'b0,x217}<<<3'd3)+$signed({1'b0,x21});
assign sharing148 = $signed({1'b0,x464})+$signed(-{1'b0,x204})+$signed(-{3'b0,x221}<<<3'd2)+$signed({2'b0,x201}<<<3'd1)+$signed(-{1'b0,x26})+$signed(-{2'b0,x439}<<<3'd1);
assign sharing149 = $signed(-{2'b0,x219}<<<3'd1)+$signed(-{1'b0,x383})+$signed({3'b0,x311}<<<3'd2)+$signed(-{2'b0,x119}<<<3'd1)+$signed(-{1'b0,x487});
assign sharing150 = $signed(-{4'b0,x408}<<<3'd3)+$signed({3'b0,x276}<<<3'd2)+$signed({2'b0,x244}<<<3'd1)+$signed(-{3'b0,x356}<<<3'd2)+$signed(-{3'b0,x485}<<<3'd2);
assign sharing151 = $signed({3'b0,x208}<<<3'd2)+$signed({2'b0,x380}<<<3'd1)+$signed(-{1'b0,x488})+$signed(-{2'b0,x297}<<<3'd1)+$signed(-{1'b0,x33})+$signed(-{1'b0,x355})+$signed({1'b0,x119});
assign sharing152 = $signed({4'b0,x452}<<<3'd3)+$signed({2'b0,x156}<<<3'd1)+$signed(-{2'b0,x44}<<<3'd1)+$signed({4'b0,x465}<<<3'd3)+$signed({3'b0,x210}<<<3'd2)+$signed(-{1'b0,x14})+$signed({1'b0,x123});
assign sharing153 = $signed(-{3'b0,x32}<<<3'd2)+$signed({1'b0,x420})+$signed({2'b0,x393}<<<3'd1)+$signed(-{1'b0,x153})+$signed(-{3'b0,x362}<<<3'd2);
assign sharing154 = $signed(-{3'b0,x244}<<<3'd2)+$signed(-{2'b0,x160}<<<3'd1)+$signed(-{2'b0,x92}<<<3'd1)+$signed(-{3'b0,x211}<<<3'd2)+$signed({1'b0,x379});
assign sharing155 = $signed(-{2'b0,x424}<<<3'd1)+$signed(-{1'b0,x208})+$signed({3'b0,x178}<<<3'd2)+$signed(-{2'b0,x314}<<<3'd1)+$signed({2'b0,x228}<<<3'd1)+$signed({2'b0,x444}<<<3'd1)+$signed({3'b0,x101}<<<3'd2)+$signed(-{3'b0,x134}<<<3'd2);
assign sharing156 = $signed(-{4'b0,x321}<<<3'd3)+$signed(-{3'b0,x70}<<<3'd2)+$signed({1'b0,x377})+$signed({3'b0,x4}<<<3'd2)+$signed({3'b0,x220}<<<3'd2)+$signed(-{3'b0,x228}<<<3'd2)+$signed(-{3'b0,x198}<<<3'd2)+$signed({3'b0,x14}<<<3'd2)+$signed(-{3'b0,x254}<<<3'd2);
assign sharing157 = $signed(-{4'b0,x460}<<<3'd3)+$signed({1'b0,x64})+$signed({1'b0,x184})+$signed({3'b0,x325}<<<3'd2)+$signed({2'b0,x493}<<<3'd1)+$signed(-{1'b0,x69})+$signed(-{3'b0,x338}<<<3'd2)+$signed(-{4'b0,x407}<<<3'd3)+$signed({3'b0,x215}<<<3'd2);
assign sharing158 = $signed(-{1'b0,x309})+$signed({3'b0,x174}<<<3'd2)+$signed({2'b0,x414}<<<3'd1)+$signed({1'b0,x270})+$signed(-{1'b0,x434});
assign sharing159 = $signed({3'b0,x478}<<<3'd2)+$signed({2'b0,x46}<<<3'd1)+$signed(-{1'b0,x388})+$signed(-{2'b0,x109}<<<3'd1);
assign sharing160 = $signed(-{4'b0,x241}<<<3'd3)+$signed({3'b0,x81}<<<3'd2)+$signed({2'b0,x43}<<<3'd1);
assign sharing161 = $signed({3'b0,x216}<<<3'd2)+$signed({1'b0,x396})+$signed({1'b0,x180})+$signed(-{3'b0,x85}<<<3'd2)+$signed(-{1'b0,x169})+$signed({2'b0,x370}<<<3'd1);
assign sharing162 = $signed({1'b0,x149})+$signed({1'b0,x493})+$signed(-{2'b0,x281}<<<3'd1)+$signed(-{3'b0,x38}<<<3'd2)+$signed({2'b0,x242}<<<3'd1)+$signed(-{3'b0,x151}<<<3'd2);
assign sharing163 = $signed(-{1'b0,x116})+$signed({3'b0,x309}<<<3'd2)+$signed({2'b0,x349}<<<3'd1)+$signed({1'b0,x369})+$signed(-{3'b0,x91}<<<3'd2);
assign sharing164 = $signed(-{3'b0,x430}<<<3'd2)+$signed(-{2'b0,x31}<<<3'd1)+$signed({2'b0,x55}<<<3'd1)+$signed(-{1'b0,x19});
assign sharing165 = $signed(-{2'b0,x176}<<<3'd1)+$signed(-{2'b0,x184}<<<3'd1)+$signed(-{2'b0,x476}<<<3'd1)+$signed(-{2'b0,x401}<<<3'd1)+$signed(-{1'b0,x385})+$signed({2'b0,x327}<<<3'd1)+$signed(-{1'b0,x427});
assign sharing166 = $signed(-{1'b0,x94})+$signed({2'b0,x110}<<<3'd1)+$signed({1'b0,x456});
assign sharing167 = $signed({3'b0,x472}<<<3'd2)+$signed({1'b0,x9})+$signed(-{1'b0,x105})+$signed(-{4'b0,x317}<<<3'd3)+$signed(-{2'b0,x29}<<<3'd1)+$signed(-{3'b0,x294}<<<3'd2)+$signed(-{2'b0,x382}<<<3'd1)+$signed({3'b0,x391}<<<3'd2);
assign sharing168 = $signed({2'b0,x328}<<<3'd1)+$signed({1'b0,x248})+$signed({3'b0,x193}<<<3'd2)+$signed({1'b0,x305})+$signed({3'b0,x52}<<<3'd2)+$signed({2'b0,x180}<<<3'd1)+$signed({2'b0,x471}<<<3'd1)+$signed({1'b0,x263});
assign sharing169 = $signed({2'b0,x352}<<<3'd1)+$signed(-{2'b0,x286}<<<3'd1)+$signed(-{1'b0,x361});
assign sharing170 = $signed({3'b0,x408}<<<3'd2)+$signed({2'b0,x208}<<<3'd1)+$signed({1'b0,x80})+$signed(-{2'b0,x266}<<<3'd1);
assign sharing171 = $signed(-{3'b0,x488}<<<3'd2)+$signed({3'b0,x113}<<<3'd2)+$signed({1'b0,x219})+$signed({2'b0,x231}<<<3'd1)+$signed({3'b0,x317}<<<3'd2)+$signed({3'b0,x413}<<<3'd2)+$signed({1'b0,x269})+$signed({3'b0,x398}<<<3'd2)+$signed({2'b0,x167}<<<3'd1);
assign sharing172 = $signed({1'b0,x8})+$signed({1'b0,x308})+$signed(-{1'b0,x140})+$signed({2'b0,x169}<<<3'd1)+$signed({2'b0,x113}<<<3'd1)+$signed({2'b0,x193}<<<3'd1)+$signed(-{1'b0,x54})+$signed({2'b0,x111}<<<3'd1);
assign sharing173 = $signed({2'b0,x168}<<<3'd1)+$signed(-{2'b0,x72}<<<3'd1)+$signed(-{1'b0,x221})+$signed({2'b0,x398}<<<3'd1)+$signed(-{4'b0,x299}<<<3'd3);
assign sharing174 = $signed({2'b0,x176}<<<3'd1)+$signed(-{1'b0,x24})+$signed({1'b0,x443});
assign sharing175 = $signed(-{3'b0,x48}<<<3'd2)+$signed({2'b0,x384}<<<3'd1)+$signed({2'b0,x143}<<<3'd1);
assign sharing176 = $signed(-{1'b0,x0})+$signed(-{1'b0,x80})+$signed({1'b0,x6})+$signed({2'b0,x481}<<<3'd1);
assign sharing177 = $signed({3'b0,x170}<<<3'd2)+$signed({2'b0,x322}<<<3'd1)+$signed(-{2'b0,x23}<<<3'd1);
assign sharing178 = $signed(-{3'b0,x195}<<<3'd2)+$signed(-{2'b0,x64}<<<3'd1)+$signed(-{1'b0,x194})+$signed(-{3'b0,x183}<<<3'd2);
assign sharing179 = $signed({3'b0,x132}<<<3'd2)+$signed(-{2'b0,x162}<<<3'd1)+$signed(-{3'b0,x140}<<<3'd2)+$signed({1'b0,x37});
assign sharing180 = $signed({2'b0,x364}<<<3'd1)+$signed({2'b0,x254}<<<3'd1)+$signed({1'b0,x420})+$signed({3'b0,x73}<<<3'd2);
assign sharing181 = $signed({3'b0,x448}<<<3'd2)+$signed({3'b0,x185}<<<3'd2)+$signed(-{3'b0,x214}<<<3'd2)+$signed({1'b0,x106})+$signed(-{4'b0,x471}<<<3'd3)+$signed(-{2'b0,x195}<<<3'd1);
assign sharing182 = $signed(-{2'b0,x0}<<<3'd1)+$signed(-{3'b0,x265}<<<3'd2)+$signed({2'b0,x238}<<<3'd1)+$signed(-{1'b0,x382})+$signed(-{2'b0,x95}<<<3'd1);
assign sharing183 = $signed({2'b0,x314}<<<3'd1)+$signed(-{3'b0,x371}<<<3'd2)+$signed(-{1'b0,x435});
assign sharing184 = $signed({1'b0,x214})+$signed(-{1'b0,x12})+$signed({3'b0,x237}<<<3'd2)+$signed({1'b0,x198})+$signed({4'b0,x255}<<<3'd3)+$signed(-{2'b0,x7}<<<3'd1)+$signed(-{1'b0,x151});
assign sharing185 = $signed(-{3'b0,x93}<<<3'd2)+$signed(-{2'b0,x469}<<<3'd1)+$signed(-{3'b0,x162}<<<3'd2)+$signed(-{1'b0,x23})+$signed({1'b0,x419});
assign sharing186 = $signed({2'b0,x66}<<<3'd1)+$signed({1'b0,x262})+$signed(-{1'b0,x203})+$signed({1'b0,x95});
assign sharing187 = $signed({4'b0,x414}<<<3'd3)+$signed(-{3'b0,x152}<<<3'd2)+$signed(-{4'b0,x205}<<<3'd3);
assign sharing188 = $signed(-{4'b0,x232}<<<3'd3)+$signed({2'b0,x76}<<<3'd1)+$signed(-{3'b0,x489}<<<3'd2)+$signed(-{3'b0,x349}<<<3'd2)+$signed(-{1'b0,x381})+$signed(-{3'b0,x427}<<<3'd2);
assign sharing189 = $signed({1'b0,x72})+$signed(-{2'b0,x389}<<<3'd1)+$signed({1'b0,x1})+$signed({2'b0,x142}<<<3'd1)+$signed({1'b0,x218})+$signed({2'b0,x139}<<<3'd1);
assign sharing190 = $signed(-{3'b0,x310}<<<3'd2)+$signed(-{2'b0,x141}<<<3'd1)+$signed(-{1'b0,x409})+$signed({4'b0,x482}<<<3'd3)+$signed(-{3'b0,x414}<<<3'd2)+$signed(-{1'b0,x293})+$signed(-{3'b0,x71}<<<3'd2);
assign sharing191 = $signed({3'b0,x192}<<<3'd2)+$signed({2'b0,x200}<<<3'd1)+$signed({1'b0,x136})+$signed(-{2'b0,x16}<<<3'd1)+$signed(-{1'b0,x215});
assign sharing192 = $signed({3'b0,x254}<<<3'd2)+$signed({4'b0,x357}<<<3'd3)+$signed(-{3'b0,x280}<<<3'd2);
assign sharing193 = $signed({3'b0,x104}<<<3'd2)+$signed(-{1'b0,x338})+$signed({3'b0,x270}<<<3'd2);
assign sharing194 = $signed(-{3'b0,x58}<<<3'd2)+$signed(-{4'b0,x161}<<<3'd3)+$signed({2'b0,x295}<<<3'd1);
assign sharing195 = $signed(-{3'b0,x96}<<<3'd2)+$signed({2'b0,x106}<<<3'd1)+$signed(-{3'b0,x477}<<<3'd2)+$signed(-{1'b0,x285});
assign sharing196 = $signed(-{2'b0,x484}<<<3'd1)+$signed({3'b0,x133}<<<3'd2)+$signed(-{1'b0,x225})+$signed(-{2'b0,x54}<<<3'd1)+$signed(-{3'b0,x107}<<<3'd2)+$signed(-{2'b0,x419}<<<3'd1);
assign sharing197 = $signed({3'b0,x50}<<<3'd2)+$signed(-{3'b0,x447}<<<3'd2)+$signed({2'b0,x337}<<<3'd1)+$signed(-{1'b0,x453});
assign sharing198 = $signed({2'b0,x108}<<<3'd1)+$signed({1'b0,x373})+$signed({2'b0,x100}<<<3'd1);
assign sharing199 = $signed({3'b0,x304}<<<3'd2)+$signed(-{1'b0,x18})+$signed({1'b0,x433});
assign sharing200 = $signed(-{2'b0,x317}<<<3'd1)+$signed({1'b0,x72})+$signed({1'b0,x436})+$signed({1'b0,x101});
assign sharing201 = $signed(-{3'b0,x332}<<<3'd2)+$signed(-{1'b0,x78})+$signed({4'b0,x7}<<<3'd3)+$signed(-{3'b0,x459}<<<3'd2)+$signed(-{1'b0,x343});
assign sharing202 = $signed(-{2'b0,x192}<<<3'd1)+$signed(-{3'b0,x157}<<<3'd2)+$signed({2'b0,x397}<<<3'd1)+$signed(-{3'b0,x171}<<<3'd2);
assign sharing203 = $signed({3'b0,x90}<<<3'd2)+$signed(-{2'b0,x285}<<<3'd1)+$signed({3'b0,x271}<<<3'd2)+$signed(-{2'b0,x307}<<<3'd1);
assign sharing204 = $signed(-{2'b0,x12}<<<3'd1)+$signed(-{1'b0,x228})+$signed(-{1'b0,x232})+$signed(-{2'b0,x284}<<<3'd1)+$signed({1'b0,x402})+$signed({1'b0,x303});
assign sharing205 = $signed({1'b0,x490})+$signed({2'b0,x235}<<<3'd1)+$signed({2'b0,x335}<<<3'd1);
assign sharing206 = $signed({2'b0,x280}<<<3'd1)+$signed({1'b0,x328})+$signed({2'b0,x274}<<<3'd1)+$signed(-{1'b0,x302})+$signed(-{3'b0,x307}<<<3'd2)+$signed(-{1'b0,x287});
assign sharing207 = $signed(-{3'b0,x421}<<<3'd2)+$signed(-{3'b0,x65}<<<3'd2)+$signed({2'b0,x57}<<<3'd1);
assign sharing208 = $signed(-{1'b0,x273})+$signed({2'b0,x197}<<<3'd1)+$signed({1'b0,x11});
assign sharing209 = $signed(-{3'b0,x305}<<<3'd2)+$signed({3'b0,x241}<<<3'd2)+$signed(-{2'b0,x269}<<<3'd1);
assign sharing210 = $signed({3'b0,x392}<<<3'd2)+$signed({2'b0,x34}<<<3'd1)+$signed({1'b0,x66})+$signed({3'b0,x159}<<<3'd2)+$signed(-{3'b0,x239}<<<3'd2);
assign sharing211 = $signed({3'b0,x236}<<<3'd2)+$signed({2'b0,x40}<<<3'd1)+$signed({1'b0,x375})+$signed({2'b0,x2}<<<3'd1)+$signed({3'b0,x203}<<<3'd2)+$signed({1'b0,x107});
assign sharing212 = $signed(-{2'b0,x318}<<<3'd1)+$signed(-{1'b0,x312})+$signed({3'b0,x231}<<<3'd2);
assign sharing213 = $signed(-{1'b0,x364})+$signed({3'b0,x83}<<<3'd2)+$signed({3'b0,x161}<<<3'd2);
assign sharing214 = $signed({3'b0,x342}<<<3'd2)+$signed({3'b0,x40}<<<3'd2)+$signed(-{3'b0,x149}<<<3'd2)+$signed({3'b0,x111}<<<3'd2);
assign sharing215 = $signed(-{3'b0,x202}<<<3'd2)+$signed({1'b0,x104})+$signed({4'b0,x291}<<<3'd3);
assign sharing216 = $signed(-{1'b0,x132})+$signed(-{1'b0,x260})+$signed({3'b0,x245}<<<3'd2)+$signed(-{3'b0,x194}<<<3'd2)+$signed({1'b0,x183});
assign sharing217 = $signed({2'b0,x470}<<<3'd1)+$signed(-{1'b0,x416})+$signed({3'b0,x387}<<<3'd2)+$signed({1'b0,x125});
assign sharing218 = $signed({2'b0,x354}<<<3'd1)+$signed({2'b0,x357}<<<3'd1)+$signed(-{2'b0,x84}<<<3'd1)+$signed({2'b0,x53}<<<3'd1);
assign sharing219 = $signed(-{2'b0,x272}<<<3'd1)+$signed({1'b0,x393})+$signed(-{3'b0,x418}<<<3'd2)+$signed({2'b0,x118}<<<3'd1)+$signed(-{2'b0,x283}<<<3'd1);
assign sharing220 = $signed(-{1'b0,x457})+$signed(-{3'b0,x277}<<<3'd2)+$signed(-{2'b0,x391}<<<3'd1)+$signed({1'b0,x275});
assign sharing221 = $signed({1'b0,x142})+$signed(-{3'b0,x416}<<<3'd2)+$signed({1'b0,x284})+$signed({1'b0,x475});
assign sharing222 = $signed({3'b0,x442}<<<3'd2)+$signed(-{2'b0,x202}<<<3'd1)+$signed(-{3'b0,x26}<<<3'd2)+$signed(-{1'b0,x237});
assign sharing223 = $signed({3'b0,x370}<<<3'd2)+$signed({3'b0,x487}<<<3'd2)+$signed(-{3'b0,x218}<<<3'd2);
assign sharing224 = $signed(-{2'b0,x65}<<<3'd1)+$signed({3'b0,x187}<<<3'd2)+$signed({2'b0,x443}<<<3'd1)+$signed({1'b0,x495});
assign sharing225 = $signed(-{3'b0,x404}<<<3'd2)+$signed({3'b0,x268}<<<3'd2)+$signed({1'b0,x168})+$signed(-{2'b0,x85}<<<3'd1);
assign sharing226 = $signed(-{2'b0,x136}<<<3'd1)+$signed(-{2'b0,x130}<<<3'd1)+$signed({2'b0,x33}<<<3'd1)+$signed(-{2'b0,x50}<<<3'd1)+$signed({2'b0,x270}<<<3'd1);
assign sharing227 = $signed({3'b0,x419}<<<3'd2)+$signed(-{1'b0,x53})+$signed(-{4'b0,x186}<<<3'd3)+$signed({3'b0,x135}<<<3'd2)+$signed(-{2'b0,x63}<<<3'd1);
assign sharing228 = $signed(-{2'b0,x368}<<<3'd1)+$signed(-{4'b0,x129}<<<3'd3)+$signed(-{1'b0,x337});
assign sharing229 = $signed(-{1'b0,x187})+$signed({2'b0,x171}<<<3'd1)+$signed({1'b0,x327});
assign sharing230 = $signed(-{3'b0,x482}<<<3'd2)+$signed({2'b0,x174}<<<3'd1)+$signed(-{1'b0,x126})+$signed({3'b0,x45}<<<3'd2);
assign sharing231 = $signed(-{4'b0,x487}<<<3'd3)+$signed({3'b0,x57}<<<3'd2)+$signed({2'b0,x213}<<<3'd1)+$signed(-{1'b0,x15});
assign sharing232 = $signed(-{1'b0,x81})+$signed(-{2'b0,x179}<<<3'd1)+$signed({1'b0,x321});
assign sharing233 = $signed({4'b0,x250}<<<3'd3)+$signed({2'b0,x360}<<<3'd1)+$signed(-{2'b0,x89}<<<3'd1);
assign sharing234 = $signed(-{4'b0,x468}<<<3'd3)+$signed(-{3'b0,x212}<<<3'd2)+$signed({2'b0,x421}<<<3'd1)+$signed(-{1'b0,x117});
assign sharing235 = $signed({3'b0,x300}<<<3'd2)+$signed(-{1'b0,x462})+$signed(-{2'b0,x251}<<<3'd1);
assign sharing236 = $signed({4'b0,x8}<<<3'd3)+$signed({1'b0,x455})+$signed(-{1'b0,x75})+$signed({1'b0,x167});
assign sharing237 = $signed(-{3'b0,x476}<<<3'd2)+$signed({2'b0,x98}<<<3'd1)+$signed(-{1'b0,x139});
assign sharing238 = $signed(-{3'b0,x145}<<<3'd2)+$signed({3'b0,x313}<<<3'd2)+$signed({2'b0,x267}<<<3'd1)+$signed(-{2'b0,x323}<<<3'd1);
assign sharing239 = $signed({4'b0,x170}<<<3'd3)+$signed({4'b0,x188}<<<3'd3)+$signed(-{3'b0,x62}<<<3'd2)+$signed({2'b0,x161}<<<3'd1);
assign sharing240 = $signed({2'b0,x132}<<<3'd1)+$signed(-{1'b0,x67})+$signed(-{2'b0,x209}<<<3'd1)+$signed({1'b0,x235});
assign sharing241 = $signed({4'b0,x116}<<<3'd3)+$signed(-{3'b0,x243}<<<3'd2)+$signed(-{1'b0,x429});
assign sharing242 = $signed({3'b0,x172}<<<3'd2)+$signed({1'b0,x404})+$signed({2'b0,x21}<<<3'd1)+$signed(-{1'b0,x5});
assign sharing243 = $signed(-{3'b0,x9}<<<3'd2)+$signed({3'b0,x55}<<<3'd2)+$signed({1'b0,x307});
assign sharing244 = $signed(-{3'b0,x376}<<<3'd2)+$signed(-{3'b0,x110}<<<3'd2)+$signed(-{4'b0,x3}<<<3'd3)+$signed(-{1'b0,x467});
assign sharing245 = $signed({2'b0,x26}<<<3'd1)+$signed({1'b0,x442})+$signed({3'b0,x415}<<<3'd2);
assign sharing246 = $signed(-{3'b0,x446}<<<3'd2)+$signed(-{1'b0,x365})+$signed(-{1'b0,x351});
assign sharing247 = $signed(-{2'b0,x298}<<<3'd1)+$signed({1'b0,x304})+$signed({1'b0,x65});
assign sharing248 = $signed(-{3'b0,x436}<<<3'd2)+$signed({2'b0,x420}<<<3'd1)+$signed({2'b0,x479}<<<3'd1);
assign sharing249 = $signed(-{4'b0,x296}<<<3'd3)+$signed({2'b0,x400}<<<3'd1)+$signed(-{3'b0,x189}<<<3'd2)+$signed({2'b0,x429}<<<3'd1);
assign sharing250 = $signed({3'b0,x177}<<<3'd2)+$signed({2'b0,x353}<<<3'd1)+$signed({2'b0,x135}<<<3'd1);
assign sharing251 = $signed({3'b0,x318}<<<3'd2)+$signed(-{3'b0,x484}<<<3'd2)+$signed({2'b0,x475}<<<3'd1);
assign sharing252 = $signed({2'b0,x58}<<<3'd1)+$signed({1'b0,x484})+$signed(-{2'b0,x36}<<<3'd1);
assign sharing253 = $signed({4'b0,x181}<<<3'd3)+$signed({3'b0,x121}<<<3'd2)+$signed({1'b0,x403});
assign sharing254 = $signed(-{3'b0,x154}<<<3'd2)+$signed({3'b0,x469}<<<3'd2)+$signed(-{1'b0,x115});
assign sharing255 = $signed({1'b0,x73})+$signed(-{1'b0,x387})+$signed({3'b0,x375}<<<3'd2)+$signed({1'b0,x25});
assign sharing256 = $signed(-{2'b0,x127}<<<3'd1)+$signed({2'b0,x297}<<<3'd1)+$signed({1'b0,x197});
assign sharing257 = $signed(-{3'b0,x148}<<<3'd2)+$signed(-{2'b0,x356}<<<3'd1)+$signed({2'b0,x371}<<<3'd1);
assign sharing258 = $signed(-{3'b0,x382}<<<3'd2)+$signed({2'b0,x287}<<<3'd1)+$signed(-{1'b0,x447});
assign sharing259 = $signed(-{3'b0,x369}<<<3'd2)+$signed({3'b0,x94}<<<3'd2)+$signed({3'b0,x89}<<<3'd2);
wire signed[14:0] temp_y  [0:19];
assign temp_y[0] = 
$signed({1'b0,x97})+$signed(-{1'b0,x322})+$signed({1'b0,x66})+$signed({3'b0,x131}<<<3'd2)+$signed({2'b0,x291}<<<3'd1)+$signed({1'b0,x3})+$signed({1'b0,x67})+$signed(-{1'b0,x292})+$signed(-{4'b0,x261}<<<3'd3)+$signed(-{4'b0,x453}<<<3'd3)+$signed(-{4'b0,x101}<<<3'd3)+$signed(-{4'b0,x134}<<<3'd3)+$signed({1'b0,x326})+$signed(-{3'b0,x392}<<<3'd2)+$signed(-{1'b0,x200})+$signed(-{4'b0,x265}<<<3'd3)+$signed(-{3'b0,x9}<<<3'd2)+$signed(-{2'b0,x169}<<<3'd1)+$signed({3'b0,x396}<<<3'd2)+$signed({1'b0,x236})+$signed(-{2'b0,x462}<<<3'd1)+$signed(-{1'b0,x175})+$signed(-{4'b0,x80}<<<3'd3)+$signed({1'b0,x112})+$signed(-{1'b0,x465})+$signed(-{3'b0,x210}<<<3'd2)+$signed({2'b0,x178}<<<3'd1)+$signed(-{3'b0,x434}<<<3'd2)+$signed(-{3'b0,x435}<<<3'd2)+$signed(-{2'b0,x339}<<<3'd1)+$signed({3'b0,x341}<<<3'd2)+$signed(-{3'b0,x309}<<<3'd2)+$signed(-{1'b0,x181})+$signed(-{4'b0,x119}<<<3'd3)+$signed(-{3'b0,x279}<<<3'd2)+$signed(-{3'b0,x247}<<<3'd2)+$signed(-{1'b0,x471})+$signed(-{3'b0,x440}<<<3'd2)+$signed({2'b0,x24}<<<3'd1)+$signed({1'b0,x122})+$signed(-{2'b0,x28}<<<3'd1)+$signed(-{1'b0,x156})+$signed(-{4'b0,x125}<<<3'd3)+$signed(-{3'b0,x317}<<<3'd2)+$signed(-{2'b0,x189}<<<3'd1)+$signed(-{3'b0,x30}<<<3'd2)+$signed({1'b0,x414})+$signed(-{4'b0,x383}<<<3'd3)+$signed(sharing8)+$signed(sharing9)+$signed(sharing36)+$signed(sharing37)+$signed(sharing50)+$signed(sharing51)+$signed(sharing66)+$signed(sharing67)+$signed(sharing90)+$signed(-sharing91)+$signed(sharing110)+$signed(sharing111)+$signed(sharing121)+$signed(sharing122)+$signed(sharing146)+$signed(sharing147)+$signed(sharing165)+$signed(sharing179)+$signed(sharing180)+$signed(sharing204)+$signed(sharing219)+$signed(sharing220)+$signed(sharing230)+$signed(sharing231)+$signed(sharing239)+$signed(sharing247)+$signed(-sharing256)+$signed(sharing258)-$signed(14'd16);
assign y0=temp_y[0][14] ==1'b1 ? 6'd0 :  
    temp_y[0][10] ==1'b1 ? 6'd63 : 
    temp_y[0][3]==1'b1 ? temp_y[0][9:4]+1'b1 : temp_y[0][9:4];
assign temp_y[1] = 
$signed(-{3'b0,x1}<<<3'd2)+$signed({1'b0,x417})+$signed({3'b0,x258}<<<3'd2)+$signed(-{2'b0,x34}<<<3'd1)+$signed({1'b0,x450})+$signed({1'b0,x259})+$signed(-{3'b0,x388}<<<3'd2)+$signed({2'b0,x260}<<<3'd1)+$signed({1'b0,x452})+$signed(-{2'b0,x5}<<<3'd1)+$signed(-{4'b0,x390}<<<3'd3)+$signed(-{2'b0,x102}<<<3'd1)+$signed(-{2'b0,x166}<<<3'd1)+$signed(-{2'b0,x8}<<<3'd1)+$signed({1'b0,x40})+$signed({1'b0,x488})+$signed({3'b0,x329}<<<3'd2)+$signed({3'b0,x233}<<<3'd2)+$signed(-{2'b0,x201}<<<3'd1)+$signed(-{4'b0,x426}<<<3'd3)+$signed(-{2'b0,x328}<<<3'd1)+$signed({1'b0,x42})+$signed({4'b0,x43}<<<3'd3)+$signed({3'b0,x235}<<<3'd2)+$signed({2'b0,x363}<<<3'd1)+$signed(-{1'b0,x138})+$signed(-{4'b0,x11}<<<3'd3)+$signed(-{1'b0,x202})+$signed({1'b0,x172})+$signed(-{3'b0,x365}<<<3'd2)+$signed({3'b0,x142}<<<3'd2)+$signed(-{2'b0,x366}<<<3'd1)+$signed({4'b0,x15}<<<3'd3)+$signed({3'b0,x399}<<<3'd2)+$signed(-{3'b0,x48}<<<3'd2)+$signed(-{3'b0,x306}<<<3'd2)+$signed({2'b0,x82}<<<3'd1)+$signed(-{2'b0,x403}<<<3'd1)+$signed({2'b0,x245}<<<3'd1)+$signed({3'b0,x22}<<<3'd2)+$signed({2'b0,x278}<<<3'd1)+$signed({2'b0,x438}<<<3'd1)+$signed(-{3'b0,x183}<<<3'd2)+$signed({1'b0,x120})+$signed(-{2'b0,x315}<<<3'd1)+$signed({3'b0,x284}<<<3'd2)+$signed(-{4'b0,x93}<<<3'd3)+$signed({3'b0,x221}<<<3'd2)+$signed({4'b0,x382}<<<3'd3)+$signed(-{3'b0,x286}<<<3'd2)+$signed({4'b0,x191}<<<3'd3)+$signed(-{3'b0,x95}<<<3'd2)+$signed(sharing14)+$signed(sharing15)+$signed(sharing22)+$signed(-sharing23)+$signed(sharing46)+$signed(sharing47)+$signed(sharing68)+$signed(sharing69)+$signed(sharing98)+$signed(-sharing99)+$signed(sharing116)+$signed(sharing117)+$signed(sharing126)+$signed(sharing127)+$signed(sharing154)+$signed(sharing155)+$signed(sharing163)+$signed(sharing164)+$signed(sharing179)+$signed(-sharing180)+$signed(sharing196)+$signed(sharing228)+$signed(sharing229)+$signed(sharing232)+$signed(sharing244)+$signed(14'd8);
assign y1=temp_y[1][14] ==1'b1 ? 6'd0 :  
    temp_y[1][10] ==1'b1 ? 6'd63 : 
    temp_y[1][3]==1'b1 ? temp_y[1][9:4]+1'b1 : temp_y[1][9:4];
assign temp_y[2] = 
$signed(-{2'b0,x160}<<<3'd1)+$signed({1'b0,x352})+$signed(-{2'b0,x96}<<<3'd1)+$signed(-{2'b0,x193}<<<3'd1)+$signed({1'b0,x99})+$signed(-{1'b0,x227})+$signed(-{2'b0,x5}<<<3'd1)+$signed(-{1'b0,x230})+$signed({1'b0,x326})+$signed({1'b0,x103})+$signed(-{4'b0,x72}<<<3'd3)+$signed(-{1'b0,x424})+$signed({3'b0,x201}<<<3'd2)+$signed(-{1'b0,x41})+$signed({3'b0,x426}<<<3'd2)+$signed({4'b0,x459}<<<3'd3)+$signed({3'b0,x235}<<<3'd2)+$signed(-{2'b0,x171}<<<3'd1)+$signed(-{2'b0,x462}<<<3'd1)+$signed({1'b0,x143})+$signed({4'b0,x433}<<<3'd3)+$signed(-{2'b0,x17}<<<3'd1)+$signed({1'b0,x465})+$signed(-{1'b0,x434})+$signed({3'b0,x467}<<<3'd2)+$signed({2'b0,x19}<<<3'd1)+$signed({2'b0,x468}<<<3'd1)+$signed({3'b0,x53}<<<3'd2)+$signed({2'b0,x181}<<<3'd1)+$signed(-{1'b0,x149})+$signed(-{1'b0,x245})+$signed(-{3'b0,x470}<<<3'd2)+$signed(-{1'b0,x29})+$signed(-{3'b0,x248}<<<3'd2)+$signed({2'b0,x120}<<<3'd1)+$signed({1'b0,x184})+$signed({2'b0,x376}<<<3'd1)+$signed(-{3'b0,x345}<<<3'd2)+$signed({2'b0,x25}<<<3'd1)+$signed(-{3'b0,x250}<<<3'd2)+$signed(-{1'b0,x186})+$signed(-{3'b0,x219}<<<3'd2)+$signed(-{2'b0,x27}<<<3'd1)+$signed({1'b0,x379})+$signed(-{3'b0,x475}<<<3'd2)+$signed(-{1'b0,x124})+$signed(-{2'b0,x157}<<<3'd1)+$signed(-{1'b0,x125})+$signed(-{1'b0,x126})+$signed(-{1'b0,x31})+$signed({2'b0,x191}<<<3'd1)+$signed(-{1'b0,x415})+$signed(sharing18)+$signed(sharing19)+$signed(sharing34)+$signed(-sharing35)+$signed(sharing58)+$signed(sharing59)+$signed(sharing64)+$signed(-sharing65)+$signed(sharing96)+$signed(sharing97)+$signed(sharing112)+$signed(sharing113)+$signed(sharing125)+$signed(sharing142)+$signed(sharing143)+$signed(sharing161)+$signed(sharing182)+$signed(-sharing183)+$signed(sharing197)+$signed(-sharing198)+$signed(sharing224)+$signed(14'd32);
assign y2=temp_y[2][14] ==1'b1 ? 6'd0 :  
    temp_y[2][10] ==1'b1 ? 6'd63 : 
    temp_y[2][3]==1'b1 ? temp_y[2][9:4]+1'b1 : temp_y[2][9:4];
assign temp_y[3] = 
$signed({1'b0,x320})+$signed(-{2'b0,x289}<<<3'd1)+$signed({2'b0,x1}<<<3'd1)+$signed({4'b0,x290}<<<3'd3)+$signed({2'b0,x226}<<<3'd1)+$signed({1'b0,x130})+$signed(-{1'b0,x195})+$signed({3'b0,x166}<<<3'd2)+$signed(-{1'b0,x198})+$signed({1'b0,x486})+$signed({3'b0,x423}<<<3'd2)+$signed({1'b0,x358})+$signed({3'b0,x39}<<<3'd2)+$signed({3'b0,x359}<<<3'd2)+$signed({1'b0,x135})+$signed({2'b0,x296}<<<3'd1)+$signed({4'b0,x329}<<<3'd3)+$signed(-{3'b0,x491}<<<3'd2)+$signed(-{1'b0,x395})+$signed({3'b0,x364}<<<3'd2)+$signed(-{2'b0,x396}<<<3'd1)+$signed({1'b0,x460})+$signed({3'b0,x173}<<<3'd2)+$signed({1'b0,x365})+$signed({1'b0,x430})+$signed({2'b0,x47}<<<3'd1)+$signed({1'b0,x79})+$signed({3'b0,x16}<<<3'd2)+$signed({1'b0,x336})+$signed(-{1'b0,x240})+$signed({3'b0,x113}<<<3'd2)+$signed({2'b0,x49}<<<3'd1)+$signed({2'b0,x177}<<<3'd1)+$signed({2'b0,x338}<<<3'd1)+$signed({4'b0,x179}<<<3'd3)+$signed(-{3'b0,x51}<<<3'd2)+$signed(-{1'b0,x19})+$signed({1'b0,x438})+$signed({3'b0,x408}<<<3'd2)+$signed({2'b0,x120}<<<3'd1)+$signed(-{2'b0,x312}<<<3'd1)+$signed(-{1'b0,x344})+$signed(-{3'b0,x153}<<<3'd2)+$signed({2'b0,x121}<<<3'd1)+$signed(-{2'b0,x25}<<<3'd1)+$signed(-{2'b0,x473}<<<3'd1)+$signed(-{3'b0,x474}<<<3'd2)+$signed({1'b0,x90})+$signed(-{1'b0,x154})+$signed({3'b0,x123}<<<3'd2)+$signed(-{2'b0,x27}<<<3'd1)+$signed(-{1'b0,x91})+$signed({3'b0,x92}<<<3'd2)+$signed(-{2'b0,x61}<<<3'd1)+$signed(-{2'b0,x255}<<<3'd1)+$signed(-{1'b0,x127})+$signed(sharing16)+$signed(-sharing17)+$signed(sharing26)+$signed(sharing27)+$signed(sharing42)+$signed(sharing43)+$signed(sharing70)+$signed(-sharing71)+$signed(sharing92)+$signed(-sharing93)+$signed(sharing110)+$signed(-sharing111)+$signed(sharing128)+$signed(sharing129)+$signed(sharing148)+$signed(-sharing149)+$signed(sharing158)+$signed(sharing176)+$signed(sharing205)+$signed(sharing206)+$signed(sharing217)+$signed(sharing218)+$signed(sharing225)+$signed(sharing233)+$signed(-sharing244)-$signed(14'd24);
assign y3=temp_y[3][14] ==1'b1 ? 6'd0 :  
    temp_y[3][10] ==1'b1 ? 6'd63 : 
    temp_y[3][3]==1'b1 ? temp_y[3][9:4]+1'b1 : temp_y[3][9:4];
assign temp_y[4] = 
$signed({4'b0,x96}<<<3'd3)+$signed({3'b0,x64}<<<3'd2)+$signed({2'b0,x480}<<<3'd1)+$signed(-{2'b0,x322}<<<3'd1)+$signed(-{1'b0,x162})+$signed(-{2'b0,x355}<<<3'd1)+$signed({3'b0,x164}<<<3'd2)+$signed({1'b0,x388})+$signed(-{1'b0,x4})+$signed(-{3'b0,x229}<<<3'd2)+$signed(-{4'b0,x102}<<<3'd3)+$signed({1'b0,x454})+$signed({4'b0,x199}<<<3'd3)+$signed(-{4'b0,x391}<<<3'd3)+$signed(-{2'b0,x359}<<<3'd1)+$signed(-{1'b0,x39})+$signed({1'b0,x103})+$signed({3'b0,x200}<<<3'd2)+$signed(-{4'b0,x9}<<<3'd3)+$signed({3'b0,x137}<<<3'd2)+$signed(-{3'b0,x265}<<<3'd2)+$signed({1'b0,x489})+$signed(-{1'b0,x425})+$signed({1'b0,x234})+$signed(-{4'b0,x268}<<<3'd3)+$signed({3'b0,x236}<<<3'd2)+$signed({1'b0,x76})+$signed(-{1'b0,x300})+$signed({3'b0,x13}<<<3'd2)+$signed(-{3'b0,x429}<<<3'd2)+$signed(-{2'b0,x77}<<<3'd1)+$signed(-{3'b0,x175}<<<3'd2)+$signed(-{2'b0,x79}<<<3'd1)+$signed({3'b0,x80}<<<3'd2)+$signed(-{3'b0,x176}<<<3'd2)+$signed(-{3'b0,x273}<<<3'd2)+$signed(-{2'b0,x241}<<<3'd1)+$signed({1'b0,x50})+$signed({3'b0,x276}<<<3'd2)+$signed({1'b0,x52})+$signed(-{3'b0,x181}<<<3'd2)+$signed({4'b0,x374}<<<3'd3)+$signed({3'b0,x150}<<<3'd2)+$signed(-{2'b0,x246}<<<3'd1)+$signed(-{1'b0,x22})+$signed({4'b0,x343}<<<3'd3)+$signed(-{3'b0,x23}<<<3'd2)+$signed(-{1'b0,x375})+$signed(-{3'b0,x248}<<<3'd2)+$signed({2'b0,x88}<<<3'd1)+$signed(-{1'b0,x472})+$signed(-{1'b0,x249})+$signed(-{4'b0,x27}<<<3'd3)+$signed(-{4'b0,x283}<<<3'd3)+$signed({2'b0,x188}<<<3'd1)+$signed({2'b0,x380}<<<3'd1)+$signed({2'b0,x381}<<<3'd1)+$signed({1'b0,x317})+$signed({2'b0,x190}<<<3'd1)+$signed(-{4'b0,x223}<<<3'd3)+$signed(-{2'b0,x447}<<<3'd1)+$signed(sharing12)+$signed(sharing13)+$signed(sharing20)+$signed(sharing21)+$signed(sharing50)+$signed(-sharing51)+$signed(sharing60)+$signed(sharing61)+$signed(sharing82)+$signed(sharing83)+$signed(sharing106)+$signed(sharing107)+$signed(sharing136)+$signed(-sharing137)+$signed(sharing154)+$signed(-sharing155)+$signed(sharing162)+$signed(sharing189)+$signed(-sharing190)+$signed(sharing202)+$signed(-sharing203)+$signed(sharing217)+$signed(-sharing218)+$signed(-sharing224)+$signed(sharing234)+$signed(sharing245)+$signed(-sharing254)+$signed(sharing257)+$signed(14'd8);
assign y4=temp_y[4][14] ==1'b1 ? 6'd0 :  
    temp_y[4][10] ==1'b1 ? 6'd63 : 
    temp_y[4][3]==1'b1 ? temp_y[4][9:4]+1'b1 : temp_y[4][9:4];
assign temp_y[5] = 
$signed(-{4'b0,x32}<<<3'd3)+$signed({3'b0,x288}<<<3'd2)+$signed({2'b0,x0}<<<3'd1)+$signed({1'b0,x96})+$signed(-{4'b0,x160}<<<3'd3)+$signed(-{2'b0,x448}<<<3'd1)+$signed(-{4'b0,x352}<<<3'd3)+$signed(-{4'b0,x225}<<<3'd3)+$signed({4'b0,x98}<<<3'd3)+$signed(-{3'b0,x129}<<<3'd2)+$signed(-{2'b0,x385}<<<3'd1)+$signed(-{3'b0,x2}<<<3'd2)+$signed(-{2'b0,x450}<<<3'd1)+$signed({3'b0,x259}<<<3'd2)+$signed({2'b0,x483}<<<3'd1)+$signed(-{3'b0,x3}<<<3'd2)+$signed(-{3'b0,x67}<<<3'd2)+$signed(-{4'b0,x68}<<<3'd3)+$signed(-{1'b0,x36})+$signed(-{4'b0,x165}<<<3'd3)+$signed(-{4'b0,x71}<<<3'd3)+$signed({2'b0,x455}<<<3'd1)+$signed(-{2'b0,x327}<<<3'd1)+$signed({3'b0,x104}<<<3'd2)+$signed({3'b0,x201}<<<3'd2)+$signed({1'b0,x170})+$signed(-{4'b0,x139}<<<3'd3)+$signed({3'b0,x363}<<<3'd2)+$signed({1'b0,x108})+$signed(-{1'b0,x205})+$signed(-{4'b0,x270}<<<3'd3)+$signed({2'b0,x206}<<<3'd1)+$signed({2'b0,x431}<<<3'd1)+$signed(-{2'b0,x16}<<<3'd1)+$signed({1'b0,x464})+$signed({4'b0,x433}<<<3'd3)+$signed(-{3'b0,x17}<<<3'd2)+$signed(-{3'b0,x465}<<<3'd2)+$signed({1'b0,x305})+$signed(-{1'b0,x146})+$signed(-{4'b0,x20}<<<3'd3)+$signed({1'b0,x468})+$signed(-{3'b0,x53}<<<3'd2)+$signed(-{3'b0,x438}<<<3'd2)+$signed({2'b0,x150}<<<3'd1)+$signed(-{1'b0,x311})+$signed({4'b0,x248}<<<3'd3)+$signed(-{4'b0,x472}<<<3'd3)+$signed({3'b0,x281}<<<3'd2)+$signed({2'b0,x442}<<<3'd1)+$signed(-{1'b0,x30})+$signed(-{4'b0,x155}<<<3'd3)+$signed(-{4'b0,x348}<<<3'd3)+$signed({2'b0,x60}<<<3'd1)+$signed(-{1'b0,x380})+$signed(-{4'b0,x350}<<<3'd3)+$signed(-{1'b0,x222})+$signed(sharing0)+$signed(-sharing1)+$signed(sharing32)+$signed(-sharing33)+$signed(sharing40)+$signed(-sharing41)+$signed(sharing60)+$signed(-sharing61)+$signed(sharing94)+$signed(sharing95)+$signed(sharing116)+$signed(-sharing117)+$signed(sharing134)+$signed(sharing135)+$signed(sharing156)+$signed(-sharing157)+$signed(sharing172)+$signed(-sharing173)+$signed(-sharing184)+$signed(sharing205)+$signed(-sharing206)+$signed(sharing216)+$signed(sharing230)+$signed(-sharing231)+$signed(sharing238)+$signed(sharing249)+$signed(-sharing253)-$signed(14'd16);
assign y5=temp_y[5][14] ==1'b1 ? 6'd0 :  
    temp_y[5][10] ==1'b1 ? 6'd63 : 
    temp_y[5][3]==1'b1 ? temp_y[5][9:4]+1'b1 : temp_y[5][9:4];
assign temp_y[6] = 
$signed({2'b0,x224}<<<3'd1)+$signed(-{2'b0,x256}<<<3'd1)+$signed({3'b0,x1}<<<3'd2)+$signed(-{2'b0,x225}<<<3'd1)+$signed({1'b0,x449})+$signed({1'b0,x353})+$signed(-{1'b0,x163})+$signed({3'b0,x255}<<<3'd2)+$signed(-{2'b0,x325}<<<3'd1)+$signed({3'b0,x326}<<<3'd2)+$signed(-{2'b0,x390}<<<3'd1)+$signed(-{1'b0,x102})+$signed(-{3'b0,x360}<<<3'd2)+$signed(-{1'b0,x233})+$signed({1'b0,x234})+$signed(-{1'b0,x202})+$signed({3'b0,x267}<<<3'd2)+$signed(-{4'b0,x75}<<<3'd3)+$signed({1'b0,x171})+$signed({3'b0,x140}<<<3'd2)+$signed({1'b0,x269})+$signed({2'b0,x366}<<<3'd1)+$signed(-{2'b0,x78}<<<3'd1)+$signed({4'b0,x111}<<<3'd3)+$signed(-{3'b0,x303}<<<3'd2)+$signed({2'b0,x207}<<<3'd1)+$signed(-{1'b0,x399})+$signed({3'b0,x336}<<<3'd2)+$signed({1'b0,x144})+$signed({1'b0,x48})+$signed(-{3'b0,x209}<<<3'd2)+$signed({2'b0,x305}<<<3'd1)+$signed({1'b0,x17})+$signed(-{2'b0,x145}<<<3'd1)+$signed({1'b0,x114})+$signed({1'b0,x370})+$signed(-{1'b0,x82})+$signed({3'b0,x180}<<<3'd2)+$signed(-{2'b0,x404}<<<3'd1)+$signed(-{1'b0,x148})+$signed(-{2'b0,x373}<<<3'd1)+$signed({1'b0,x342})+$signed(-{1'b0,x61})+$signed({1'b0,x215})+$signed({4'b0,x376}<<<3'd3)+$signed({1'b0,x93})+$signed(-{2'b0,x24}<<<3'd1)+$signed({3'b0,x441}<<<3'd2)+$signed(-{3'b0,x186}<<<3'd2)+$signed({1'b0,x314})+$signed({4'b0,x123}<<<3'd3)+$signed(-{1'b0,x250})+$signed(-{1'b0,x189})+$signed(-{3'b0,x155}<<<3'd2)+$signed(-{3'b0,x347}<<<3'd2)+$signed({2'b0,x476}<<<3'd1)+$signed(-{1'b0,x316})+$signed({3'b0,x381}<<<3'd2)+$signed(-{2'b0,x253}<<<3'd1)+$signed(-{1'b0,x445})+$signed(-{4'b0,x446}<<<3'd3)+$signed({1'b0,x414})+$signed({3'b0,x31}<<<3'd2)+$signed(sharing4)+$signed(-sharing5)+$signed(sharing26)+$signed(-sharing27)+$signed(sharing52)+$signed(-sharing53)+$signed(sharing74)+$signed(-sharing75)+$signed(sharing84)+$signed(-sharing85)+$signed(sharing112)+$signed(-sharing113)+$signed(sharing134)+$signed(-sharing135)+$signed(sharing150)+$signed(-sharing151)+$signed(sharing159)+$signed(-sharing160)+$signed(sharing177)+$signed(-sharing178)+$signed(sharing199)+$signed(-sharing200)+$signed(sharing210)+$signed(sharing221)+$signed(-sharing234)+$signed(sharing243)+$signed(sharing252)-$signed(14'd48);
assign y6=temp_y[6][14] ==1'b1 ? 6'd0 :  
    temp_y[6][10] ==1'b1 ? 6'd63 : 
    temp_y[6][3]==1'b1 ? temp_y[6][9:4]+1'b1 : temp_y[6][9:4];
assign temp_y[7] = 
$signed({3'b0,x320}<<<3'd2)+$signed({4'b0,x385}<<<3'd3)+$signed({3'b0,x321}<<<3'd2)+$signed({2'b0,x225}<<<3'd1)+$signed({1'b0,x418})+$signed({1'b0,x482})+$signed(-{2'b0,x3}<<<3'd1)+$signed({3'b0,x420}<<<3'd2)+$signed(-{3'b0,x292}<<<3'd2)+$signed(-{3'b0,x228}<<<3'd2)+$signed(-{1'b0,x485})+$signed(-{1'b0,x325})+$signed({2'b0,x134}<<<3'd1)+$signed(-{3'b0,x327}<<<3'd2)+$signed(-{4'b0,x488}<<<3'd3)+$signed(-{4'b0,x201}<<<3'd3)+$signed({3'b0,x393}<<<3'd2)+$signed(-{2'b0,x457}<<<3'd1)+$signed({1'b0,x297})+$signed(-{2'b0,x489}<<<3'd1)+$signed({2'b0,x42}<<<3'd1)+$signed({2'b0,x234}<<<3'd1)+$signed(-{2'b0,x138}<<<3'd1)+$signed({1'b0,x395})+$signed({4'b0,x460}<<<3'd3)+$signed({4'b0,x333}<<<3'd3)+$signed(-{2'b0,x109}<<<3'd1)+$signed({2'b0,x430}<<<3'd1)+$signed(-{1'b0,x366})+$signed(-{4'b0,x303}<<<3'd3)+$signed(-{2'b0,x271}<<<3'd1)+$signed(-{3'b0,x112}<<<3'd2)+$signed(-{4'b0,x305}<<<3'd3)+$signed(-{3'b0,x401}<<<3'd2)+$signed({2'b0,x306}<<<3'd1)+$signed(-{2'b0,x434}<<<3'd1)+$signed(-{4'b0,x403}<<<3'd3)+$signed(-{4'b0,x435}<<<3'd3)+$signed(-{3'b0,x20}<<<3'd2)+$signed({2'b0,x276}<<<3'd1)+$signed(-{1'b0,x308})+$signed({2'b0,x149}<<<3'd1)+$signed({2'b0,x277}<<<3'd1)+$signed({1'b0,x54})+$signed({2'b0,x87}<<<3'd1)+$signed({1'b0,x441})+$signed({1'b0,x158})+$signed({3'b0,x122}<<<3'd2)+$signed(-{2'b0,x91}<<<3'd1)+$signed(-{2'b0,x59}<<<3'd1)+$signed(-{2'b0,x379}<<<3'd1)+$signed({3'b0,x156}<<<3'd2)+$signed({1'b0,x60})+$signed({1'b0,x380})+$signed(-{3'b0,x349}<<<3'd2)+$signed(-{4'b0,x414}<<<3'd3)+$signed({1'b0,x222})+$signed({1'b0,x287})+$signed(sharing14)+$signed(-sharing15)+$signed(sharing20)+$signed(-sharing21)+$signed(sharing54)+$signed(-sharing55)+$signed(sharing66)+$signed(-sharing67)+$signed(sharing80)+$signed(-sharing81)+$signed(sharing102)+$signed(-sharing103)+$signed(sharing130)+$signed(-sharing131)+$signed(sharing142)+$signed(-sharing143)+$signed(sharing166)+$signed(-sharing167)+$signed(sharing185)+$signed(-sharing186)+$signed(sharing201)+$signed(sharing216)+$signed(-sharing222)+$signed(sharing233)+$signed(sharing246)+$signed(sharing252)+$signed(14'd16);
assign y7=temp_y[7][14] ==1'b1 ? 6'd0 :  
    temp_y[7][10] ==1'b1 ? 6'd63 : 
    temp_y[7][3]==1'b1 ? temp_y[7][9:4]+1'b1 : temp_y[7][9:4];
assign temp_y[8] = 
$signed({4'b0,x320}<<<3'd3)+$signed(-{4'b0,x224}<<<3'd3)+$signed({2'b0,x288}<<<3'd1)+$signed({1'b0,x192})+$signed({2'b0,x416}<<<3'd1)+$signed({2'b0,x386}<<<3'd1)+$signed({2'b0,x418}<<<3'd1)+$signed({3'b0,x3}<<<3'd2)+$signed({4'b0,x4}<<<3'd3)+$signed({4'b0,x292}<<<3'd3)+$signed(-{1'b0,x452})+$signed({3'b0,x165}<<<3'd2)+$signed(-{3'b0,x453}<<<3'd2)+$signed({4'b0,x70}<<<3'd3)+$signed(-{2'b0,x454}<<<3'd1)+$signed({3'b0,x199}<<<3'd2)+$signed({3'b0,x71}<<<3'd2)+$signed({1'b0,x489})+$signed(-{1'b0,x297})+$signed(-{1'b0,x10})+$signed(-{1'b0,x170})+$signed(-{3'b0,x75}<<<3'd2)+$signed(-{4'b0,x491}<<<3'd3)+$signed(-{1'b0,x299})+$signed(-{4'b0,x492}<<<3'd3)+$signed({4'b0,x45}<<<3'd3)+$signed({2'b0,x173}<<<3'd1)+$signed(-{1'b0,x301})+$signed({1'b0,x367})+$signed(-{2'b0,x432}<<<3'd1)+$signed({4'b0,x337}<<<3'd3)+$signed(-{4'b0,x242}<<<3'd3)+$signed({4'b0,x339}<<<3'd3)+$signed({3'b0,x211}<<<3'd2)+$signed(-{4'b0,x243}<<<3'd3)+$signed(-{2'b0,x275}<<<3'd1)+$signed({4'b0,x84}<<<3'd3)+$signed({2'b0,x372}<<<3'd1)+$signed({3'b0,x85}<<<3'd2)+$signed({2'b0,x309}<<<3'd1)+$signed(-{4'b0,x278}<<<3'd3)+$signed({3'b0,x22}<<<3'd2)+$signed({2'b0,x214}<<<3'd1)+$signed(-{4'b0,x310}<<<3'd3)+$signed(-{1'b0,x374})+$signed({1'b0,x183})+$signed(-{3'b0,x282}<<<3'd2)+$signed(-{3'b0,x122}<<<3'd2)+$signed({3'b0,x315}<<<3'd2)+$signed({2'b0,x188}<<<3'd1)+$signed({1'b0,x220})+$signed({2'b0,x252}<<<3'd1)+$signed({4'b0,x253}<<<3'd3)+$signed(-{3'b0,x29}<<<3'd2)+$signed(-{2'b0,x285}<<<3'd1)+$signed({3'b0,x63}<<<3'd2)+$signed(-{3'b0,x479}<<<3'd2)+$signed(-{1'b0,x349})+$signed(sharing10)+$signed(sharing11)+$signed(sharing30)+$signed(sharing31)+$signed(sharing44)+$signed(sharing45)+$signed(sharing62)+$signed(sharing63)+$signed(sharing90)+$signed(sharing91)+$signed(sharing114)+$signed(sharing115)+$signed(sharing132)+$signed(sharing133)+$signed(sharing148)+$signed(sharing149)+$signed(sharing168)+$signed(sharing169)+$signed(sharing182)+$signed(sharing183)+$signed(sharing199)+$signed(sharing200)+$signed(sharing214)+$signed(sharing215)+$signed(sharing226)+$signed(sharing235)+$signed(sharing249)+$signed(sharing254)+$signed(sharing259)+$signed(14'd24);
assign y8=temp_y[8][14] ==1'b1 ? 6'd0 :  
    temp_y[8][10] ==1'b1 ? 6'd63 : 
    temp_y[8][3]==1'b1 ? temp_y[8][9:4]+1'b1 : temp_y[8][9:4];
assign temp_y[9] = 
$signed(-{4'b0,x448}<<<3'd3)+$signed(-{3'b0,x352}<<<3'd2)+$signed(-{2'b0,x480}<<<3'd1)+$signed(-{4'b0,x97}<<<3'd3)+$signed({3'b0,x225}<<<3'd2)+$signed(-{2'b0,x449}<<<3'd1)+$signed(-{2'b0,x417}<<<3'd1)+$signed(-{4'b0,x450}<<<3'd3)+$signed(-{3'b0,x66}<<<3'd2)+$signed({3'b0,x386}<<<3'd2)+$signed(-{3'b0,x322}<<<3'd2)+$signed({3'b0,x354}<<<3'd2)+$signed({3'b0,x451}<<<3'd2)+$signed({1'b0,x259})+$signed(-{4'b0,x324}<<<3'd3)+$signed({2'b0,x228}<<<3'd1)+$signed(-{1'b0,x68})+$signed({1'b0,x389})+$signed({1'b0,x325})+$signed(-{2'b0,x262}<<<3'd1)+$signed(-{4'b0,x359}<<<3'd3)+$signed({1'b0,x391})+$signed(-{4'b0,x200}<<<3'd3)+$signed(-{3'b0,x328}<<<3'd2)+$signed(-{3'b0,x424}<<<3'd2)+$signed(-{3'b0,x393}<<<3'd2)+$signed({3'b0,x266}<<<3'd2)+$signed(-{4'b0,x267}<<<3'd3)+$signed(-{4'b0,x363}<<<3'd3)+$signed({3'b0,x492}<<<3'd2)+$signed(-{4'b0,x461}<<<3'd3)+$signed({3'b0,x397}<<<3'd2)+$signed(-{3'b0,x205}<<<3'd2)+$signed({1'b0,x13})+$signed({2'b0,x237}<<<3'd1)+$signed(-{3'b0,x334}<<<3'd2)+$signed(-{2'b0,x14}<<<3'd1)+$signed(-{1'b0,x206})+$signed(-{4'b0,x302}<<<3'd3)+$signed({3'b0,x494}<<<3'd2)+$signed({1'b0,x431})+$signed(-{4'b0,x16}<<<3'd3)+$signed(-{4'b0,x272}<<<3'd3)+$signed(-{1'b0,x47})+$signed(-{1'b0,x432})+$signed(-{2'b0,x17}<<<3'd1)+$signed({4'b0,x50}<<<3'd3)+$signed({3'b0,x18}<<<3'd2)+$signed(-{4'b0,x51}<<<3'd3)+$signed(-{3'b0,x339}<<<3'd2)+$signed(-{4'b0,x307}<<<3'd3)+$signed({1'b0,x83})+$signed(-{4'b0,x180}<<<3'd3)+$signed(-{3'b0,x308}<<<3'd2)+$signed(-{4'b0,x244}<<<3'd3)+$signed(-{4'b0,x213}<<<3'd3)+$signed({3'b0,x309}<<<3'd2)+$signed(-{2'b0,x341}<<<3'd1)+$signed({3'b0,x279}<<<3'd2)+$signed(-{3'b0,x439}<<<3'd2)+$signed({1'b0,x407})+$signed({3'b0,x248}<<<3'd2)+$signed(-{4'b0,x409}<<<3'd3)+$signed(-{4'b0,x442}<<<3'd3)+$signed({1'b0,x282})+$signed(-{4'b0,x315}<<<3'd3)+$signed(-{3'b0,x126}<<<3'd2)+$signed({2'b0,x94}<<<3'd1)+$signed({3'b0,x284}<<<3'd2)+$signed({2'b0,x220}<<<3'd1)+$signed(-{2'b0,x477}<<<3'd1)+$signed(-{1'b0,x413})+$signed({3'b0,x350}<<<3'd2)+$signed({2'b0,x478}<<<3'd1)+$signed(sharing0)+$signed(sharing1)+$signed(sharing24)+$signed(sharing25)+$signed(sharing48)+$signed(sharing49)+$signed(sharing70)+$signed(sharing71)+$signed(sharing84)+$signed(sharing85)+$signed(sharing108)+$signed(sharing109)+$signed(sharing132)+$signed(-sharing133)+$signed(sharing144)+$signed(-sharing145)+$signed(sharing162)+$signed(sharing174)+$signed(sharing175)+$signed(sharing201)+$signed(sharing208)+$signed(sharing209)+$signed(sharing223)+$signed(sharing236)+$signed(sharing247)+$signed(14'd8);
assign y9=temp_y[9][14] ==1'b1 ? 6'd0 :  
    temp_y[9][10] ==1'b1 ? 6'd63 : 
    temp_y[9][3]==1'b1 ? temp_y[9][9:4]+1'b1 : temp_y[9][9:4];
assign temp_y[10] = 
$signed(-{1'b0,x160})+$signed({3'b0,x481}<<<3'd2)+$signed({2'b0,x2}<<<3'd1)+$signed(-{3'b0,x323}<<<3'd2)+$signed({2'b0,x259}<<<3'd1)+$signed(-{3'b0,x293}<<<3'd2)+$signed({3'b0,x6}<<<3'd2)+$signed(-{2'b0,x38}<<<3'd1)+$signed({2'b0,x166}<<<3'd1)+$signed({2'b0,x487}<<<3'd1)+$signed({3'b0,x8}<<<3'd2)+$signed({1'b0,x137})+$signed({1'b0,x201})+$signed(-{2'b0,x330}<<<3'd1)+$signed(-{1'b0,x298})+$signed(-{2'b0,x395}<<<3'd1)+$signed(-{1'b0,x107})+$signed(-{2'b0,x460}<<<3'd1)+$signed(-{1'b0,x268})+$signed(-{3'b0,x301}<<<3'd2)+$signed({2'b0,x461}<<<3'd1)+$signed({3'b0,x430}<<<3'd2)+$signed({3'b0,x78}<<<3'd2)+$signed({3'b0,x206}<<<3'd2)+$signed({1'b0,x110})+$signed(-{1'b0,x463})+$signed({2'b0,x304}<<<3'd1)+$signed({1'b0,x208})+$signed(-{2'b0,x210}<<<3'd1)+$signed(-{2'b0,x466}<<<3'd1)+$signed(-{3'b0,x211}<<<3'd2)+$signed(-{3'b0,x371}<<<3'd2)+$signed(-{3'b0,x84}<<<3'd2)+$signed({2'b0,x405}<<<3'd1)+$signed({1'b0,x277})+$signed({4'b0,x342}<<<3'd3)+$signed(-{2'b0,x311}<<<3'd1)+$signed({1'b0,x247})+$signed(-{3'b0,x120}<<<3'd2)+$signed({3'b0,x409}<<<3'd2)+$signed(-{2'b0,x441}<<<3'd1)+$signed(-{1'b0,x313})+$signed(-{1'b0,x121})+$signed({2'b0,x314}<<<3'd1)+$signed({1'b0,x474})+$signed({3'b0,x251}<<<3'd2)+$signed(-{3'b0,x27}<<<3'd2)+$signed(-{2'b0,x156}<<<3'd1)+$signed(-{2'b0,x124}<<<3'd1)+$signed({3'b0,x253}<<<3'd2)+$signed(-{2'b0,x221}<<<3'd1)+$signed({3'b0,x478}<<<3'd2)+$signed(-{2'b0,x446}<<<3'd1)+$signed(-{2'b0,x159}<<<3'd1)+$signed(sharing16)+$signed(sharing17)+$signed(sharing32)+$signed(sharing33)+$signed(sharing48)+$signed(-sharing49)+$signed(sharing76)+$signed(-sharing77)+$signed(sharing80)+$signed(sharing81)+$signed(sharing104)+$signed(-sharing105)+$signed(sharing121)+$signed(-sharing122)+$signed(sharing138)+$signed(sharing139)+$signed(sharing161)+$signed(sharing177)+$signed(sharing178)+$signed(sharing202)+$signed(sharing203)+$signed(sharing212)+$signed(sharing213)+$signed(sharing232)+$signed(sharing241)+$signed(sharing255)+$signed(sharing259)+$signed(14'd56);
assign y10=temp_y[10][14] ==1'b1 ? 6'd0 :  
    temp_y[10][10] ==1'b1 ? 6'd63 : 
    temp_y[10][3]==1'b1 ? temp_y[10][9:4]+1'b1 : temp_y[10][9:4];
assign temp_y[11] = 
$signed(-{4'b0,x96}<<<3'd3)+$signed(-{3'b0,x0}<<<3'd2)+$signed({2'b0,x97}<<<3'd1)+$signed({1'b0,x289})+$signed({1'b0,x162})+$signed({4'b0,x163}<<<3'd3)+$signed({3'b0,x388}<<<3'd2)+$signed({3'b0,x295}<<<3'd2)+$signed(-{1'b0,x7})+$signed({1'b0,x359})+$signed(-{1'b0,x296})+$signed({3'b0,x457}<<<3'd2)+$signed({2'b0,x9}<<<3'd1)+$signed(-{1'b0,x201})+$signed(-{1'b0,x329})+$signed(-{1'b0,x330})+$signed(-{1'b0,x43})+$signed(-{3'b0,x12}<<<3'd2)+$signed({1'b0,x268})+$signed({2'b0,x301}<<<3'd1)+$signed({1'b0,x173})+$signed({1'b0,x493})+$signed({3'b0,x78}<<<3'd2)+$signed({1'b0,x334})+$signed({3'b0,x207}<<<3'd2)+$signed({2'b0,x15}<<<3'd1)+$signed({2'b0,x336}<<<3'd1)+$signed({2'b0,x241}<<<3'd1)+$signed(-{1'b0,x49})+$signed(-{4'b0,x114}<<<3'd3)+$signed({3'b0,x275}<<<3'd2)+$signed({2'b0,x467}<<<3'd1)+$signed({3'b0,x115}<<<3'd2)+$signed(-{3'b0,x244}<<<3'd2)+$signed({2'b0,x340}<<<3'd1)+$signed({1'b0,x277})+$signed({1'b0,x85})+$signed({1'b0,x469})+$signed({3'b0,x118}<<<3'd2)+$signed(-{2'b0,x279}<<<3'd1)+$signed(-{2'b0,x215}<<<3'd1)+$signed({2'b0,x442}<<<3'd1)+$signed({1'b0,x27})+$signed({3'b0,x348}<<<3'd2)+$signed(-{3'b0,x252}<<<3'd2)+$signed({1'b0,x476})+$signed({1'b0,x188})+$signed(sharing18)+$signed(-sharing19)+$signed(sharing38)+$signed(sharing39)+$signed(sharing42)+$signed(-sharing43)+$signed(sharing74)+$signed(sharing75)+$signed(sharing86)+$signed(sharing87)+$signed(sharing102)+$signed(sharing103)+$signed(sharing120)+$signed(sharing152)+$signed(sharing153)+$signed(sharing168)+$signed(-sharing169)+$signed(sharing174)+$signed(-sharing175)+$signed(sharing192)+$signed(-sharing193)+$signed(sharing211)+$signed(sharing227)+$signed(-sharing240)+$signed(sharing253)+$signed(-sharing258)-$signed(14'd48);
assign y11=temp_y[11][14] ==1'b1 ? 6'd0 :  
    temp_y[11][10] ==1'b1 ? 6'd63 : 
    temp_y[11][3]==1'b1 ? temp_y[11][9:4]+1'b1 : temp_y[11][9:4];
assign temp_y[12] = 
$signed({2'b0,x128}<<<3'd1)+$signed({1'b0,x64})+$signed(-{1'b0,x224})+$signed({3'b0,x417}<<<3'd2)+$signed({3'b0,x34}<<<3'd2)+$signed({3'b0,x482}<<<3'd2)+$signed(-{3'b0,x99}<<<3'd2)+$signed(-{2'b0,x483}<<<3'd1)+$signed(-{4'b0,x100}<<<3'd3)+$signed({2'b0,x388}<<<3'd1)+$signed({1'b0,x350})+$signed(-{2'b0,x485}<<<3'd1)+$signed(-{3'b0,x488}<<<3'd2)+$signed({3'b0,x361}<<<3'd2)+$signed(-{4'b0,x362}<<<3'd3)+$signed({2'b0,x234}<<<3'd1)+$signed({1'b0,x298})+$signed(-{2'b0,x490}<<<3'd1)+$signed({1'b0,x267})+$signed({1'b0,x108})+$signed({4'b0,x173}<<<3'd3)+$signed({1'b0,x45})+$signed({4'b0,x238}<<<3'd3)+$signed({1'b0,x46})+$signed(-{1'b0,x366})+$signed({3'b0,x143}<<<3'd2)+$signed(-{2'b0,x111}<<<3'd1)+$signed(-{1'b0,x207})+$signed({2'b0,x304}<<<3'd1)+$signed({1'b0,x16})+$signed({2'b0,x433}<<<3'd1)+$signed({1'b0,x145})+$signed({1'b0,x401})+$signed({3'b0,x146}<<<3'd2)+$signed({2'b0,x274}<<<3'd1)+$signed({4'b0,x370}<<<3'd3)+$signed(-{2'b0,x210}<<<3'd1)+$signed(-{1'b0,x306})+$signed(-{2'b0,x211}<<<3'd1)+$signed({2'b0,x308}<<<3'd1)+$signed(-{1'b0,x20})+$signed(-{1'b0,x276})+$signed(-{2'b0,x85}<<<3'd1)+$signed(-{3'b0,x406}<<<3'd2)+$signed({2'b0,x182}<<<3'd1)+$signed({2'b0,x374}<<<3'd1)+$signed(-{3'b0,x375}<<<3'd2)+$signed({2'b0,x216}<<<3'd1)+$signed({1'b0,x152})+$signed(-{2'b0,x248}<<<3'd1)+$signed({3'b0,x217}<<<3'd2)+$signed(-{3'b0,x410}<<<3'd2)+$signed({2'b0,x186}<<<3'd1)+$signed({2'b0,x187}<<<3'd1)+$signed({1'b0,x347})+$signed(-{1'b0,x219})+$signed({2'b0,x316}<<<3'd1)+$signed({1'b0,x348})+$signed(-{2'b0,x412}<<<3'd1)+$signed({3'b0,x317}<<<3'd2)+$signed(-{1'b0,x60})+$signed(-{4'b0,x189}<<<3'd3)+$signed({1'b0,x446})+$signed({2'b0,x383}<<<3'd1)+$signed(sharing4)+$signed(sharing5)+$signed(sharing38)+$signed(-sharing39)+$signed(sharing58)+$signed(-sharing59)+$signed(sharing62)+$signed(-sharing63)+$signed(sharing82)+$signed(-sharing83)+$signed(sharing100)+$signed(sharing101)+$signed(sharing123)+$signed(-sharing124)+$signed(sharing140)+$signed(sharing141)+$signed(sharing163)+$signed(-sharing164)+$signed(-sharing176)+$signed(sharing204)+$signed(sharing208)+$signed(-sharing209)+$signed(-sharing237)+$signed(sharing248)+$signed(sharing251)-$signed(14'd8);
assign y12=temp_y[12][14] ==1'b1 ? 6'd0 :  
    temp_y[12][10] ==1'b1 ? 6'd63 : 
    temp_y[12][3]==1'b1 ? temp_y[12][9:4]+1'b1 : temp_y[12][9:4];
assign temp_y[13] = 
$signed({2'b0,x96}<<<3'd1)+$signed(-{3'b0,x322}<<<3'd2)+$signed({3'b0,x66}<<<3'd2)+$signed({3'b0,x226}<<<3'd2)+$signed(-{3'b0,x130}<<<3'd2)+$signed({3'b0,x291}<<<3'd2)+$signed({3'b0,x483}<<<3'd2)+$signed(-{1'b0,x323})+$signed({3'b0,x196}<<<3'd2)+$signed({3'b0,x324}<<<3'd2)+$signed({1'b0,x100})+$signed({3'b0,x325}<<<3'd2)+$signed({2'b0,x165}<<<3'd1)+$signed(-{1'b0,x453})+$signed(-{2'b0,x133}<<<3'd1)+$signed(-{2'b0,x6}<<<3'd1)+$signed({3'b0,x199}<<<3'd2)+$signed({2'b0,x232}<<<3'd1)+$signed(-{1'b0,x8})+$signed({2'b0,x137}<<<3'd1)+$signed({2'b0,x265}<<<3'd1)+$signed({2'b0,x233}<<<3'd1)+$signed({3'b0,x138}<<<3'd2)+$signed(-{2'b0,x10}<<<3'd1)+$signed(-{4'b0,x331}<<<3'd3)+$signed({3'b0,x11}<<<3'd2)+$signed({2'b0,x459}<<<3'd1)+$signed(-{1'b0,x363})+$signed(-{3'b0,x268}<<<3'd2)+$signed({2'b0,x332}<<<3'd1)+$signed(-{2'b0,x236}<<<3'd1)+$signed({2'b0,x205}<<<3'd1)+$signed({2'b0,x365}<<<3'd1)+$signed({4'b0,x366}<<<3'd3)+$signed({3'b0,x14}<<<3'd2)+$signed({3'b0,x46}<<<3'd2)+$signed({1'b0,x494})+$signed({2'b0,x431}<<<3'd1)+$signed({1'b0,x176})+$signed({2'b0,x273}<<<3'd1)+$signed(-{2'b0,x18}<<<3'd1)+$signed(-{2'b0,x275}<<<3'd1)+$signed({1'b0,x147})+$signed(-{1'b0,x339})+$signed(-{3'b0,x52}<<<3'd2)+$signed({2'b0,x341}<<<3'd1)+$signed({1'b0,x213})+$signed(-{1'b0,x245})+$signed({3'b0,x470}<<<3'd2)+$signed({3'b0,x54}<<<3'd2)+$signed({1'b0,x86})+$signed(-{3'b0,x182}<<<3'd2)+$signed({3'b0,x343}<<<3'd2)+$signed({3'b0,x311}<<<3'd2)+$signed(-{1'b0,x150})+$signed(-{3'b0,x471}<<<3'd2)+$signed({2'b0,x153}<<<3'd1)+$signed({2'b0,x217}<<<3'd1)+$signed({3'b0,x314}<<<3'd2)+$signed({2'b0,x218}<<<3'd1)+$signed({1'b0,x378})+$signed(-{1'b0,x346})+$signed(-{3'b0,x188}<<<3'd2)+$signed(-{2'b0,x477}<<<3'd1)+$signed(-{2'b0,x445}<<<3'd1)+$signed({3'b0,x190}<<<3'd2)+$signed(-{1'b0,x62})+$signed({1'b0,x63})+$signed(sharing12)+$signed(-sharing13)+$signed(sharing36)+$signed(-sharing37)+$signed(sharing54)+$signed(sharing55)+$signed(sharing68)+$signed(-sharing69)+$signed(sharing88)+$signed(-sharing89)+$signed(sharing100)+$signed(-sharing101)+$signed(sharing120)+$signed(sharing138)+$signed(-sharing139)+$signed(sharing158)+$signed(sharing184)+$signed(sharing191)+$signed(-sharing207)+$signed(sharing221)+$signed(-sharing235)+$signed(sharing242)-$signed(14'd8);
assign y13=temp_y[13][14] ==1'b1 ? 6'd0 :  
    temp_y[13][10] ==1'b1 ? 6'd63 : 
    temp_y[13][3]==1'b1 ? temp_y[13][9:4]+1'b1 : temp_y[13][9:4];
assign temp_y[14] = 
$signed(-{4'b0,x416}<<<3'd3)+$signed({1'b0,x384})+$signed(-{1'b0,x258})+$signed(-{4'b0,x99}<<<3'd3)+$signed({3'b0,x355}<<<3'd2)+$signed(-{3'b0,x291}<<<3'd2)+$signed({1'b0,x356})+$signed(-{1'b0,x196})+$signed({3'b0,x389}<<<3'd2)+$signed(-{3'b0,x287}<<<3'd2)+$signed({4'b0,x486}<<<3'd3)+$signed({3'b0,x454}<<<3'd2)+$signed({2'b0,x230}<<<3'd1)+$signed(-{4'b0,x262}<<<3'd3)+$signed({3'b0,x327}<<<3'd2)+$signed({2'b0,x263}<<<3'd1)+$signed({1'b0,x71})+$signed(-{3'b0,x8}<<<3'd2)+$signed(-{4'b0,x169}<<<3'd3)+$signed({2'b0,x265}<<<3'd1)+$signed({2'b0,x329}<<<3'd1)+$signed({4'b0,x490}<<<3'd3)+$signed(-{3'b0,x298}<<<3'd2)+$signed({2'b0,x10}<<<3'd1)+$signed(-{3'b0,x426}<<<3'd2)+$signed({2'b0,x491}<<<3'd1)+$signed(-{1'b0,x331})+$signed({4'b0,x364}<<<3'd3)+$signed({3'b0,x204}<<<3'd2)+$signed({2'b0,x492}<<<3'd1)+$signed(-{2'b0,x140}<<<3'd1)+$signed(-{1'b0,x332})+$signed({3'b0,x493}<<<3'd2)+$signed({1'b0,x45})+$signed({2'b0,x110}<<<3'd1)+$signed(-{2'b0,x47}<<<3'd1)+$signed({3'b0,x272}<<<3'd2)+$signed(-{4'b0,x273}<<<3'd3)+$signed({3'b0,x401}<<<3'd2)+$signed({4'b0,x434}<<<3'd3)+$signed({1'b0,x274})+$signed({1'b0,x402})+$signed({4'b0,x467}<<<3'd3)+$signed({2'b0,x243}<<<3'd1)+$signed(-{3'b0,x340}<<<3'd2)+$signed({1'b0,x437})+$signed(-{1'b0,x405})+$signed({2'b0,x342}<<<3'd1)+$signed({2'b0,x182}<<<3'd1)+$signed(-{4'b0,x183}<<<3'd3)+$signed(-{4'b0,x439}<<<3'd3)+$signed(-{2'b0,x343}<<<3'd1)+$signed(-{3'b0,x217}<<<3'd2)+$signed({4'b0,x218}<<<3'd3)+$signed({3'b0,x186}<<<3'd2)+$signed(-{4'b0,x187}<<<3'd3)+$signed(-{4'b0,x251}<<<3'd3)+$signed({4'b0,x476}<<<3'd3)+$signed(-{3'b0,x380}<<<3'd2)+$signed({2'b0,x28}<<<3'd1)+$signed({4'b0,x445}<<<3'd3)+$signed({3'b0,x285}<<<3'd2)+$signed(-{3'b0,x319}<<<3'd2)+$signed(sharing6)+$signed(-sharing7)+$signed(sharing24)+$signed(-sharing25)+$signed(sharing44)+$signed(-sharing45)+$signed(sharing78)+$signed(sharing79)+$signed(sharing94)+$signed(-sharing95)+$signed(sharing106)+$signed(-sharing107)+$signed(sharing125)+$signed(sharing152)+$signed(-sharing153)+$signed(sharing170)+$signed(-sharing171)+$signed(sharing187)+$signed(-sharing188)+$signed(sharing196)+$signed(sharing210)+$signed(sharing225)+$signed(sharing239)+$signed(sharing246)+$signed(sharing255)-$signed(14'd8);
assign y14=temp_y[14][14] ==1'b1 ? 6'd0 :  
    temp_y[14][10] ==1'b1 ? 6'd63 : 
    temp_y[14][3]==1'b1 ? temp_y[14][9:4]+1'b1 : temp_y[14][9:4];
assign temp_y[15] = 
$signed({3'b0,x384}<<<3'd2)+$signed({2'b0,x320}<<<3'd1)+$signed(-{2'b0,x1}<<<3'd1)+$signed(-{1'b0,x193})+$signed(-{2'b0,x194}<<<3'd1)+$signed(-{2'b0,x290}<<<3'd1)+$signed({2'b0,x159}<<<3'd1)+$signed({2'b0,x355}<<<3'd1)+$signed(-{2'b0,x229}<<<3'd1)+$signed(-{1'b0,x133})+$signed({3'b0,x70}<<<3'd2)+$signed({1'b0,x294})+$signed({3'b0,x263}<<<3'd2)+$signed({2'b0,x103}<<<3'd1)+$signed(-{3'b0,x296}<<<3'd2)+$signed(-{2'b0,x392}<<<3'd1)+$signed({3'b0,x425}<<<3'd2)+$signed({2'b0,x41}<<<3'd1)+$signed({3'b0,x42}<<<3'd2)+$signed({3'b0,x170}<<<3'd2)+$signed({3'b0,x267}<<<3'd2)+$signed({3'b0,x363}<<<3'd2)+$signed(-{3'b0,x331}<<<3'd2)+$signed(-{3'b0,x491}<<<3'd2)+$signed(-{3'b0,x461}<<<3'd2)+$signed({2'b0,x493}<<<3'd1)+$signed(-{2'b0,x13}<<<3'd1)+$signed(-{1'b0,x109})+$signed(-{1'b0,x238})+$signed(-{4'b0,x80}<<<3'd3)+$signed(-{4'b0,x48}<<<3'd3)+$signed(-{2'b0,x240}<<<3'd1)+$signed(-{1'b0,x432})+$signed(-{4'b0,x305}<<<3'd3)+$signed(-{4'b0,x113}<<<3'd3)+$signed(-{4'b0,x369}<<<3'd3)+$signed(-{1'b0,x241})+$signed(-{3'b0,x338}<<<3'd2)+$signed(-{3'b0,x19}<<<3'd2)+$signed(-{2'b0,x339}<<<3'd1)+$signed({4'b0,x149}<<<3'd3)+$signed({2'b0,x21}<<<3'd1)+$signed(-{2'b0,x53}<<<3'd1)+$signed(-{2'b0,x437}<<<3'd1)+$signed({2'b0,x86}<<<3'd1)+$signed({1'b0,x470})+$signed({2'b0,x408}<<<3'd1)+$signed({3'b0,x281}<<<3'd2)+$signed({3'b0,x473}<<<3'd2)+$signed(-{3'b0,x377}<<<3'd2)+$signed({1'b0,x314})+$signed({4'b0,x347}<<<3'd3)+$signed(-{1'b0,x250})+$signed(-{4'b0,x30}<<<3'd3)+$signed(-{1'b0,x286})+$signed(-{4'b0,x95}<<<3'd3)+$signed(-{2'b0,x255}<<<3'd1)+$signed({1'b0,x190})+$signed(sharing10)+$signed(-sharing11)+$signed(sharing28)+$signed(-sharing29)+$signed(sharing56)+$signed(-sharing57)+$signed(sharing78)+$signed(-sharing79)+$signed(sharing96)+$signed(-sharing97)+$signed(sharing118)+$signed(-sharing119)+$signed(sharing126)+$signed(-sharing127)+$signed(sharing140)+$signed(-sharing141)+$signed(-sharing165)+$signed(-sharing181)+$signed(-sharing191)+$signed(sharing211)+$signed(sharing222)+$signed(-sharing236)+$signed(sharing241)+$signed(sharing257)+$signed(14'd56);
assign y15=temp_y[15][14] ==1'b1 ? 6'd0 :  
    temp_y[15][10] ==1'b1 ? 6'd63 : 
    temp_y[15][3]==1'b1 ? temp_y[15][9:4]+1'b1 : temp_y[15][9:4];
assign temp_y[16] = 
$signed(-{2'b0,x352}<<<3'd1)+$signed({3'b0,x385}<<<3'd2)+$signed(-{2'b0,x321}<<<3'd1)+$signed(-{1'b0,x2})+$signed(-{4'b0,x355}<<<3'd3)+$signed(-{2'b0,x35}<<<3'd1)+$signed({4'b0,x452}<<<3'd3)+$signed(-{3'b0,x68}<<<3'd2)+$signed(-{4'b0,x325}<<<3'd3)+$signed({3'b0,x37}<<<3'd2)+$signed({1'b0,x38})+$signed(-{4'b0,x135}<<<3'd3)+$signed({3'b0,x455}<<<3'd2)+$signed(-{1'b0,x296})+$signed({3'b0,x105}<<<3'd2)+$signed({2'b0,x73}<<<3'd1)+$signed({2'b0,x361}<<<3'd1)+$signed({4'b0,x138}<<<3'd3)+$signed(-{2'b0,x458}<<<3'd1)+$signed({2'b0,x427}<<<3'd1)+$signed(-{3'b0,x460}<<<3'd2)+$signed({4'b0,x494}<<<3'd3)+$signed({3'b0,x174}<<<3'd2)+$signed({3'b0,x79}<<<3'd2)+$signed({2'b0,x495}<<<3'd1)+$signed({2'b0,x463}<<<3'd1)+$signed(-{2'b0,x175}<<<3'd1)+$signed(-{1'b0,x16})+$signed(-{1'b0,x272})+$signed(-{4'b0,x466}<<<3'd3)+$signed({2'b0,x146}<<<3'd1)+$signed({1'b0,x82})+$signed({2'b0,x52}<<<3'd1)+$signed({1'b0,x84})+$signed({2'b0,x180}<<<3'd1)+$signed({4'b0,x118}<<<3'd3)+$signed({4'b0,x311}<<<3'd3)+$signed(-{1'b0,x216})+$signed(-{4'b0,x89}<<<3'd3)+$signed(-{3'b0,x153}<<<3'd2)+$signed(-{1'b0,x248})+$signed({1'b0,x28})+$signed(-{4'b0,x221}<<<3'd3)+$signed(-{2'b0,x93}<<<3'd1)+$signed({1'b0,x157})+$signed({4'b0,x158}<<<3'd3)+$signed({1'b0,x478})+$signed(-{4'b0,x63}<<<3'd3)+$signed(-{3'b0,x351}<<<3'd2)+$signed({1'b0,x349})+$signed(sharing2)+$signed(sharing3)+$signed(sharing34)+$signed(sharing35)+$signed(sharing40)+$signed(sharing41)+$signed(sharing76)+$signed(sharing77)+$signed(sharing98)+$signed(sharing99)+$signed(sharing118)+$signed(sharing119)+$signed(sharing130)+$signed(sharing131)+$signed(sharing144)+$signed(sharing145)+$signed(sharing170)+$signed(sharing171)+$signed(sharing189)+$signed(sharing190)+$signed(sharing194)+$signed(sharing195)+$signed(sharing207)+$signed(sharing226)+$signed(sharing240)+$signed(sharing243)+$signed(sharing251)+$signed(sharing256)-$signed(14'd0);
assign y16=temp_y[16][14] ==1'b1 ? 6'd0 :  
    temp_y[16][10] ==1'b1 ? 6'd63 : 
    temp_y[16][3]==1'b1 ? temp_y[16][9:4]+1'b1 : temp_y[16][9:4];
assign temp_y[17] = 
$signed(-{3'b0,x256}<<<3'd2)+$signed({3'b0,x32}<<<3'd2)+$signed({3'b0,x289}<<<3'd2)+$signed(-{2'b0,x129}<<<3'd1)+$signed({3'b0,x163}<<<3'd2)+$signed({2'b0,x99}<<<3'd1)+$signed({3'b0,x68}<<<3'd2)+$signed({2'b0,x388}<<<3'd1)+$signed({1'b0,x196})+$signed({3'b0,x357}<<<3'd2)+$signed({3'b0,x102}<<<3'd2)+$signed({1'b0,x231})+$signed(-{4'b0,x415}<<<3'd3)+$signed(-{3'b0,x264}<<<3'd2)+$signed(-{4'b0,x168}<<<3'd3)+$signed(-{3'b0,x232}<<<3'd2)+$signed({2'b0,x488}<<<3'd1)+$signed(-{3'b0,x169}<<<3'd2)+$signed(-{4'b0,x330}<<<3'd3)+$signed(-{3'b0,x266}<<<3'd2)+$signed(-{4'b0,x458}<<<3'd3)+$signed(-{4'b0,x42}<<<3'd3)+$signed(-{4'b0,x427}<<<3'd3)+$signed(-{2'b0,x11}<<<3'd1)+$signed({1'b0,x267})+$signed(-{4'b0,x396}<<<3'd3)+$signed(-{4'b0,x204}<<<3'd3)+$signed({4'b0,x364}<<<3'd3)+$signed(-{3'b0,x492}<<<3'd2)+$signed(-{1'b0,x428})+$signed({1'b0,x77})+$signed({4'b0,x495}<<<3'd3)+$signed({3'b0,x335}<<<3'd2)+$signed(-{2'b0,x399}<<<3'd1)+$signed({2'b0,x175}<<<3'd1)+$signed({4'b0,x144}<<<3'd3)+$signed(-{4'b0,x240}<<<3'd3)+$signed(-{2'b0,x208}<<<3'd1)+$signed({1'b0,x272})+$signed(-{2'b0,x464}<<<3'd1)+$signed(-{4'b0,x369}<<<3'd3)+$signed(-{2'b0,x81}<<<3'd1)+$signed({3'b0,x241}<<<3'd2)+$signed({2'b0,x114}<<<3'd1)+$signed(-{4'b0,x467}<<<3'd3)+$signed(-{3'b0,x275}<<<3'd2)+$signed(-{4'b0,x52}<<<3'd3)+$signed({3'b0,x116}<<<3'd2)+$signed(-{4'b0,x308}<<<3'd3)+$signed({4'b0,x54}<<<3'd3)+$signed(-{4'b0,x438}<<<3'd3)+$signed({2'b0,x22}<<<3'd1)+$signed(-{4'b0,x183}<<<3'd3)+$signed({3'b0,x87}<<<3'd2)+$signed(-{4'b0,x247}<<<3'd3)+$signed(-{3'b0,x119}<<<3'd2)+$signed({3'b0,x24}<<<3'd2)+$signed(-{1'b0,x376})+$signed({4'b0,x314}<<<3'd3)+$signed(-{4'b0,x379}<<<3'd3)+$signed({3'b0,x443}<<<3'd2)+$signed(-{3'b0,x60}<<<3'd2)+$signed(-{1'b0,x412})+$signed(-{4'b0,x285}<<<3'd3)+$signed({2'b0,x125}<<<3'd1)+$signed(-{4'b0,x478}<<<3'd3)+$signed({4'b0,x351}<<<3'd3)+$signed(-{1'b0,x255})+$signed(sharing8)+$signed(-sharing9)+$signed(sharing22)+$signed(sharing23)+$signed(sharing52)+$signed(sharing53)+$signed(sharing72)+$signed(sharing73)+$signed(sharing92)+$signed(sharing93)+$signed(sharing104)+$signed(sharing105)+$signed(sharing136)+$signed(sharing137)+$signed(sharing156)+$signed(sharing157)+$signed(sharing166)+$signed(sharing167)+$signed(sharing181)+$signed(sharing197)+$signed(sharing198)+$signed(sharing214)+$signed(-sharing215)+$signed(sharing227)+$signed(sharing237)+$signed(sharing242)-$signed(14'd8);
assign y17=temp_y[17][14] ==1'b1 ? 6'd0 :  
    temp_y[17][10] ==1'b1 ? 6'd63 : 
    temp_y[17][3]==1'b1 ? temp_y[17][9:4]+1'b1 : temp_y[17][9:4];
assign temp_y[18] = 
$signed(-{1'b0,x32})+$signed(-{4'b0,x417}<<<3'd3)+$signed({4'b0,x386}<<<3'd3)+$signed(-{4'b0,x418}<<<3'd3)+$signed({2'b0,x258}<<<3'd1)+$signed(-{2'b0,x66}<<<3'd1)+$signed({3'b0,x162}<<<3'd2)+$signed({3'b0,x67}<<<3'd2)+$signed({3'b0,x451}<<<3'd2)+$signed({1'b0,x131})+$signed(-{2'b0,x387}<<<3'd1)+$signed(-{2'b0,x350}<<<3'd1)+$signed({2'b0,x68}<<<3'd1)+$signed(-{1'b0,x290})+$signed(-{4'b0,x197}<<<3'd3)+$signed(-{1'b0,x35})+$signed(-{4'b0,x484}<<<3'd3)+$signed(-{4'b0,x421}<<<3'd3)+$signed(-{4'b0,x166}<<<3'd3)+$signed(-{3'b0,x198}<<<3'd2)+$signed(-{4'b0,x455}<<<3'd3)+$signed({3'b0,x136}<<<3'd2)+$signed(-{4'b0,x41}<<<3'd3)+$signed(-{3'b0,x106}<<<3'd2)+$signed({2'b0,x138}<<<3'd1)+$signed({1'b0,x362})+$signed(-{4'b0,x203}<<<3'd3)+$signed(-{2'b0,x75}<<<3'd1)+$signed({2'b0,x235}<<<3'd1)+$signed(-{3'b0,x191}<<<3'd2)+$signed({3'b0,x428}<<<3'd2)+$signed({2'b0,x300}<<<3'd1)+$signed(-{1'b0,x140})+$signed(-{4'b0,x493}<<<3'd3)+$signed({2'b0,x77}<<<3'd1)+$signed({1'b0,x397})+$signed({1'b0,x13})+$signed({4'b0,x398}<<<3'd3)+$signed({2'b0,x45}<<<3'd1)+$signed(-{1'b0,x111})+$signed({4'b0,x208}<<<3'd3)+$signed({4'b0,x176}<<<3'd3)+$signed({2'b0,x369}<<<3'd1)+$signed(-{1'b0,x209})+$signed(-{3'b0,x274}<<<3'd2)+$signed({2'b0,x402}<<<3'd1)+$signed({1'b0,x210})+$signed({1'b0,x466})+$signed(-{3'b0,x82}<<<3'd2)+$signed(-{1'b0,x178})+$signed(-{2'b0,x307}<<<3'd1)+$signed({4'b0,x212}<<<3'd3)+$signed({3'b0,x372}<<<3'd2)+$signed(-{4'b0,x277}<<<3'd3)+$signed(-{1'b0,x226})+$signed(-{4'b0,x309}<<<3'd3)+$signed({4'b0,x182}<<<3'd3)+$signed(-{4'b0,x343}<<<3'd3)+$signed({3'b0,x87}<<<3'd2)+$signed(-{4'b0,x377}<<<3'd3)+$signed(-{2'b0,x281}<<<3'd1)+$signed(-{2'b0,x89}<<<3'd1)+$signed({4'b0,x90}<<<3'd3)+$signed(-{2'b0,x474}<<<3'd1)+$signed({1'b0,x410})+$signed(-{2'b0,x347}<<<3'd1)+$signed({2'b0,x59}<<<3'd1)+$signed({4'b0,x28}<<<3'd3)+$signed({4'b0,x284}<<<3'd3)+$signed(-{4'b0,x156}<<<3'd3)+$signed({3'b0,x93}<<<3'd2)+$signed(-{3'b0,x157}<<<3'd2)+$signed({1'b0,x477})+$signed(-{4'b0,x190}<<<3'd3)+$signed(-{2'b0,x30}<<<3'd1)+$signed(-{3'b0,x127}<<<3'd2)+$signed(-{1'b0,x319})+$signed(sharing2)+$signed(-sharing3)+$signed(sharing28)+$signed(sharing29)+$signed(sharing46)+$signed(-sharing47)+$signed(sharing64)+$signed(sharing65)+$signed(sharing88)+$signed(sharing89)+$signed(sharing114)+$signed(-sharing115)+$signed(sharing123)+$signed(sharing124)+$signed(sharing146)+$signed(-sharing147)+$signed(sharing159)+$signed(sharing160)+$signed(sharing187)+$signed(sharing188)+$signed(sharing192)+$signed(sharing193)+$signed(sharing212)+$signed(-sharing213)+$signed(-sharing223)+$signed(sharing238)+$signed(sharing245)+$signed(sharing250)-$signed(14'd8);
assign y18=temp_y[18][14] ==1'b1 ? 6'd0 :  
    temp_y[18][10] ==1'b1 ? 6'd63 : 
    temp_y[18][3]==1'b1 ? temp_y[18][9:4]+1'b1 : temp_y[18][9:4];
assign temp_y[19] = 
$signed(-{4'b0,x0}<<<3'd3)+$signed(-{2'b0,x32}<<<3'd1)+$signed({1'b0,x256})+$signed(-{1'b0,x352})+$signed(-{2'b0,x160}<<<3'd1)+$signed({3'b0,x226}<<<3'd2)+$signed({1'b0,x290})+$signed({1'b0,x98})+$signed({3'b0,x101}<<<3'd2)+$signed(-{3'b0,x230}<<<3'd2)+$signed(-{1'b0,x134})+$signed(-{2'b0,x199}<<<3'd1)+$signed(-{4'b0,x73}<<<3'd3)+$signed(-{1'b0,x137})+$signed(-{1'b0,x265})+$signed({2'b0,x170}<<<3'd1)+$signed({2'b0,x268}<<<3'd1)+$signed({2'b0,x204}<<<3'd1)+$signed({1'b0,x492})+$signed(-{4'b0,x109}<<<3'd3)+$signed(-{3'b0,x269}<<<3'd2)+$signed(-{2'b0,x141}<<<3'd1)+$signed(-{4'b0,x237}<<<3'd3)+$signed({3'b0,x240}<<<3'd2)+$signed({2'b0,x80}<<<3'd1)+$signed({1'b0,x400})+$signed(-{1'b0,x176})+$signed({1'b0,x242})+$signed(-{4'b0,x19}<<<3'd3)+$signed(-{3'b0,x147}<<<3'd2)+$signed({2'b0,x51}<<<3'd1)+$signed({1'b0,x179})+$signed(-{1'b0,x211})+$signed(-{1'b0,x116})+$signed(-{2'b0,x117}<<<3'd1)+$signed({3'b0,x406}<<<3'd2)+$signed({2'b0,x310}<<<3'd1)+$signed(-{3'b0,x470}<<<3'd2)+$signed(-{1'b0,x182})+$signed(-{2'b0,x407}<<<3'd1)+$signed(-{2'b0,x375}<<<3'd1)+$signed(-{3'b0,x216}<<<3'd2)+$signed(-{3'b0,x56}<<<3'd2)+$signed(-{1'b0,x88})+$signed({1'b0,x249})+$signed(-{2'b0,x26}<<<3'd1)+$signed(-{2'b0,x378}<<<3'd1)+$signed(-{4'b0,x219}<<<3'd3)+$signed(-{3'b0,x27}<<<3'd2)+$signed({2'b0,x443}<<<3'd1)+$signed(-{3'b0,x91}<<<3'd2)+$signed(-{1'b0,x411})+$signed({3'b0,x412}<<<3'd2)+$signed({2'b0,x284}<<<3'd1)+$signed({1'b0,x124})+$signed(-{3'b0,x251}<<<3'd2)+$signed(-{1'b0,x315})+$signed({1'b0,x62})+$signed(-{1'b0,x446})+$signed({1'b0,x63})+$signed(sharing6)+$signed(sharing7)+$signed(sharing30)+$signed(-sharing31)+$signed(sharing56)+$signed(sharing57)+$signed(sharing72)+$signed(-sharing73)+$signed(sharing86)+$signed(-sharing87)+$signed(sharing108)+$signed(-sharing109)+$signed(sharing128)+$signed(-sharing129)+$signed(sharing150)+$signed(sharing151)+$signed(sharing172)+$signed(sharing173)+$signed(sharing185)+$signed(sharing186)+$signed(sharing194)+$signed(-sharing195)+$signed(sharing219)+$signed(-sharing220)+$signed(sharing228)+$signed(-sharing229)+$signed(sharing248)+$signed(sharing250)+$signed(14'd72);
assign y19=temp_y[19][14] ==1'b1 ? 6'd0 :  
    temp_y[19][10] ==1'b1 ? 6'd63 : 
    temp_y[19][3]==1'b1 ? temp_y[19][9:4]+1'b1 : temp_y[19][9:4];
endmodule