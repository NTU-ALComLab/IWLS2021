module Bind(
input [7:0] x0 ,
input [7:0] x1 ,
input [7:0] x2 ,
input [7:0] x3 ,
input [7:0] x4 ,
input [7:0] x5 ,
input [7:0] x6 ,
input [7:0] x7 ,
input [7:0] x8 ,
input [7:0] x9 ,
input [7:0] x10 ,
input [7:0] x11 ,
input [7:0] x12 ,
input [7:0] x13 ,
input [7:0] x14 ,
input [7:0] x15 ,
input [7:0] x16 ,
input [7:0] x17 ,
input [7:0] x18 ,
input [7:0] x19 ,
input [7:0] x20 ,
input [7:0] x21 ,
input [7:0] x22 ,
input [7:0] x23 ,
input [7:0] x24 ,
input [7:0] x25 ,
input [7:0] x26 ,
input [7:0] x27 ,
input [7:0] x28 ,
input [7:0] x29 ,
input [7:0] x30 ,
input [7:0] x31 ,
input [7:0] x32 ,
input [7:0] x33 ,
input [7:0] x34 ,
input [7:0] x35 ,
input [7:0] x36 ,
input [7:0] x37 ,
input [7:0] x38 ,
input [7:0] x39 ,
input [7:0] x40 ,
input [7:0] x41 ,
input [7:0] x42 ,
input [7:0] x43 ,
input [7:0] x44 ,
input [7:0] x45 ,
input [7:0] x46 ,
input [7:0] x47 ,
input [7:0] x48 ,
input [7:0] x49 ,
input [7:0] x50 ,
input [7:0] x51 ,
input [7:0] x52 ,
input [7:0] x53 ,
input [7:0] x54 ,
input [7:0] x55 ,
input [7:0] x56 ,
input [7:0] x57 ,
input [7:0] x58 ,
input [7:0] x59 ,
input [7:0] x60 ,
input [7:0] x61 ,
input [7:0] x62 ,
input [7:0] x63 ,
input [7:0] x64 ,
input [7:0] x65 ,
input [7:0] x66 ,
input [7:0] x67 ,
input [7:0] x68 ,
input [7:0] x69 ,
input [7:0] x70 ,
input [7:0] x71 ,
input [7:0] x72 ,
input [7:0] x73 ,
input [7:0] x74 ,
input [7:0] x75 ,
input [7:0] x76 ,
input [7:0] x77 ,
input [7:0] x78 ,
input [7:0] x79 ,
input [7:0] x80 ,
input [7:0] x81 ,
input [7:0] x82 ,
input [7:0] x83 ,
input [7:0] x84 ,
input [7:0] x85 ,
input [7:0] x86 ,
input [7:0] x87 ,
input [7:0] x88 ,
input [7:0] x89 ,
input [7:0] x90 ,
input [7:0] x91 ,
input [7:0] x92 ,
input [7:0] x93 ,
input [7:0] x94 ,
input [7:0] x95 ,
input [7:0] x96 ,
input [7:0] x97 ,
input [7:0] x98 ,
input [7:0] x99 ,
input [7:0] x100 ,
input [7:0] x101 ,
input [7:0] x102 ,
input [7:0] x103 ,
input [7:0] x104 ,
input [7:0] x105 ,
input [7:0] x106 ,
input [7:0] x107 ,
input [7:0] x108 ,
input [7:0] x109 ,
input [7:0] x110 ,
input [7:0] x111 ,
input [7:0] x112 ,
input [7:0] x113 ,
input [7:0] x114 ,
input [7:0] x115 ,
input [7:0] x116 ,
input [7:0] x117 ,
input [7:0] x118 ,
input [7:0] x119 ,
input [7:0] x120 ,
input [7:0] x121 ,
input [7:0] x122 ,
input [7:0] x123 ,
input [7:0] x124 ,
input [7:0] x125 ,
input [7:0] x126 ,
input [7:0] x127 ,
input [7:0] x128 ,
input [7:0] x129 ,
input [7:0] x130 ,
input [7:0] x131 ,
input [7:0] x132 ,
input [7:0] x133 ,
input [7:0] x134 ,
input [7:0] x135 ,
input [7:0] x136 ,
input [7:0] x137 ,
input [7:0] x138 ,
input [7:0] x139 ,
input [7:0] x140 ,
input [7:0] x141 ,
input [7:0] x142 ,
input [7:0] x143 ,
input [7:0] x144 ,
input [7:0] x145 ,
input [7:0] x146 ,
input [7:0] x147 ,
input [7:0] x148 ,
input [7:0] x149 ,
input [7:0] x150 ,
input [7:0] x151 ,
input [7:0] x152 ,
input [7:0] x153 ,
input [7:0] x154 ,
input [7:0] x155 ,
input [7:0] x156 ,
input [7:0] x157 ,
input [7:0] x158 ,
input [7:0] x159 ,
input [7:0] x160 ,
input [7:0] x161 ,
input [7:0] x162 ,
input [7:0] x163 ,
input [7:0] x164 ,
input [7:0] x165 ,
input [7:0] x166 ,
input [7:0] x167 ,
input [7:0] x168 ,
input [7:0] x169 ,
input [7:0] x170 ,
input [7:0] x171 ,
input [7:0] x172 ,
input [7:0] x173 ,
input [7:0] x174 ,
input [7:0] x175 ,
input [7:0] x176 ,
input [7:0] x177 ,
input [7:0] x178 ,
input [7:0] x179 ,
input [7:0] x180 ,
input [7:0] x181 ,
input [7:0] x182 ,
input [7:0] x183 ,
input [7:0] x184 ,
input [7:0] x185 ,
input [7:0] x186 ,
input [7:0] x187 ,
input [7:0] x188 ,
input [7:0] x189 ,
input [7:0] x190 ,
input [7:0] x191 ,
input [7:0] x192 ,
input [7:0] x193 ,
input [7:0] x194 ,
input [7:0] x195 ,
input [7:0] x196 ,
input [7:0] x197 ,
input [7:0] x198 ,
input [7:0] x199 ,
input [7:0] x200 ,
input [7:0] x201 ,
input [7:0] x202 ,
input [7:0] x203 ,
input [7:0] x204 ,
input [7:0] x205 ,
input [7:0] x206 ,
input [7:0] x207 ,
input [7:0] x208 ,
input [7:0] x209 ,
input [7:0] x210 ,
input [7:0] x211 ,
input [7:0] x212 ,
input [7:0] x213 ,
input [7:0] x214 ,
input [7:0] x215 ,
input [7:0] x216 ,
input [7:0] x217 ,
input [7:0] x218 ,
input [7:0] x219 ,
input [7:0] x220 ,
input [7:0] x221 ,
input [7:0] x222 ,
input [7:0] x223 ,
input [7:0] x224 ,
input [7:0] x225 ,
input [7:0] x226 ,
input [7:0] x227 ,
input [7:0] x228 ,
input [7:0] x229 ,
input [7:0] x230 ,
input [7:0] x231 ,
input [7:0] x232 ,
input [7:0] x233 ,
input [7:0] x234 ,
input [7:0] x235 ,
input [7:0] x236 ,
input [7:0] x237 ,
input [7:0] x238 ,
input [7:0] x239 ,
input [7:0] x240 ,
input [7:0] x241 ,
input [7:0] x242 ,
input [7:0] x243 ,
input [7:0] x244 ,
input [7:0] x245 ,
input [7:0] x246 ,
input [7:0] x247 ,
input [7:0] x248 ,
input [7:0] x249 ,
input [7:0] x250 ,
input [7:0] x251 ,
input [7:0] x252 ,
input [7:0] x253 ,
input [7:0] x254 ,
input [7:0] x255 ,
input [7:0] x256 ,
input [7:0] x257 ,
input [7:0] x258 ,
input [7:0] x259 ,
input [7:0] x260 ,
input [7:0] x261 ,
input [7:0] x262 ,
input [7:0] x263 ,
input [7:0] x264 ,
input [7:0] x265 ,
input [7:0] x266 ,
input [7:0] x267 ,
input [7:0] x268 ,
input [7:0] x269 ,
input [7:0] x270 ,
input [7:0] x271 ,
input [7:0] x272 ,
input [7:0] x273 ,
input [7:0] x274 ,
input [7:0] x275 ,
input [7:0] x276 ,
input [7:0] x277 ,
input [7:0] x278 ,
input [7:0] x279 ,
input [7:0] x280 ,
input [7:0] x281 ,
input [7:0] x282 ,
input [7:0] x283 ,
input [7:0] x284 ,
input [7:0] x285 ,
input [7:0] x286 ,
input [7:0] x287 ,
input [7:0] x288 ,
input [7:0] x289 ,
input [7:0] x290 ,
input [7:0] x291 ,
input [7:0] x292 ,
input [7:0] x293 ,
input [7:0] x294 ,
input [7:0] x295 ,
input [7:0] x296 ,
input [7:0] x297 ,
input [7:0] x298 ,
input [7:0] x299 ,
input [7:0] x300 ,
input [7:0] x301 ,
input [7:0] x302 ,
input [7:0] x303 ,
input [7:0] x304 ,
input [7:0] x305 ,
input [7:0] x306 ,
input [7:0] x307 ,
input [7:0] x308 ,
input [7:0] x309 ,
input [7:0] x310 ,
input [7:0] x311 ,
input [7:0] x312 ,
input [7:0] x313 ,
input [7:0] x314 ,
input [7:0] x315 ,
input [7:0] x316 ,
input [7:0] x317 ,
input [7:0] x318 ,
input [7:0] x319 ,
input [7:0] x320 ,
input [7:0] x321 ,
input [7:0] x322 ,
input [7:0] x323 ,
input [7:0] x324 ,
input [7:0] x325 ,
input [7:0] x326 ,
input [7:0] x327 ,
input [7:0] x328 ,
input [7:0] x329 ,
input [7:0] x330 ,
input [7:0] x331 ,
input [7:0] x332 ,
input [7:0] x333 ,
input [7:0] x334 ,
input [7:0] x335 ,
input [7:0] x336 ,
input [7:0] x337 ,
input [7:0] x338 ,
input [7:0] x339 ,
input [7:0] x340 ,
input [7:0] x341 ,
input [7:0] x342 ,
input [7:0] x343 ,
input [7:0] x344 ,
input [7:0] x345 ,
input [7:0] x346 ,
input [7:0] x347 ,
input [7:0] x348 ,
input [7:0] x349 ,
input [7:0] x350 ,
input [7:0] x351 ,
input [7:0] x352 ,
input [7:0] x353 ,
input [7:0] x354 ,
input [7:0] x355 ,
input [7:0] x356 ,
input [7:0] x357 ,
input [7:0] x358 ,
input [7:0] x359 ,
input [7:0] x360 ,
input [7:0] x361 ,
input [7:0] x362 ,
input [7:0] x363 ,
input [7:0] x364 ,
input [7:0] x365 ,
input [7:0] x366 ,
input [7:0] x367 ,
input [7:0] x368 ,
input [7:0] x369 ,
input [7:0] x370 ,
input [7:0] x371 ,
input [7:0] x372 ,
input [7:0] x373 ,
input [7:0] x374 ,
input [7:0] x375 ,
input [7:0] x376 ,
input [7:0] x377 ,
input [7:0] x378 ,
input [7:0] x379 ,
input [7:0] x380 ,
input [7:0] x381 ,
input [7:0] x382 ,
input [7:0] x383 ,
input [7:0] x384 ,
input [7:0] x385 ,
input [7:0] x386 ,
input [7:0] x387 ,
input [7:0] x388 ,
input [7:0] x389 ,
input [7:0] x390 ,
input [7:0] x391 ,
input [7:0] x392 ,
input [7:0] x393 ,
input [7:0] x394 ,
input [7:0] x395 ,
input [7:0] x396 ,
input [7:0] x397 ,
input [7:0] x398 ,
input [7:0] x399 ,
input [7:0] x400 ,
input [7:0] x401 ,
input [7:0] x402 ,
input [7:0] x403 ,
input [7:0] x404 ,
input [7:0] x405 ,
input [7:0] x406 ,
input [7:0] x407 ,
input [7:0] x408 ,
input [7:0] x409 ,
input [7:0] x410 ,
input [7:0] x411 ,
input [7:0] x412 ,
input [7:0] x413 ,
input [7:0] x414 ,
input [7:0] x415 ,
input [7:0] x416 ,
input [7:0] x417 ,
input [7:0] x418 ,
input [7:0] x419 ,
input [7:0] x420 ,
input [7:0] x421 ,
input [7:0] x422 ,
input [7:0] x423 ,
input [7:0] x424 ,
input [7:0] x425 ,
input [7:0] x426 ,
input [7:0] x427 ,
input [7:0] x428 ,
input [7:0] x429 ,
input [7:0] x430 ,
input [7:0] x431 ,
input [7:0] x432 ,
input [7:0] x433 ,
input [7:0] x434 ,
input [7:0] x435 ,
input [7:0] x436 ,
input [7:0] x437 ,
input [7:0] x438 ,
input [7:0] x439 ,
input [7:0] x440 ,
input [7:0] x441 ,
input [7:0] x442 ,
input [7:0] x443 ,
input [7:0] x444 ,
input [7:0] x445 ,
input [7:0] x446 ,
input [7:0] x447 ,
input [7:0] x448 ,
input [7:0] x449 ,
input [7:0] x450 ,
input [7:0] x451 ,
input [7:0] x452 ,
input [7:0] x453 ,
input [7:0] x454 ,
input [7:0] x455 ,
input [7:0] x456 ,
input [7:0] x457 ,
input [7:0] x458 ,
input [7:0] x459 ,
input [7:0] x460 ,
input [7:0] x461 ,
input [7:0] x462 ,
input [7:0] x463 ,
input [7:0] x464 ,
input [7:0] x465 ,
input [7:0] x466 ,
input [7:0] x467 ,
input [7:0] x468 ,
input [7:0] x469 ,
input [7:0] x470 ,
input [7:0] x471 ,
input [7:0] x472 ,
input [7:0] x473 ,
input [7:0] x474 ,
input [7:0] x475 ,
input [7:0] x476 ,
input [7:0] x477 ,
input [7:0] x478 ,
input [7:0] x479 ,
input [7:0] x480 ,
input [7:0] x481 ,
input [7:0] x482 ,
input [7:0] x483 ,
input [7:0] x484 ,
input [7:0] x485 ,
input [7:0] x486 ,
input [7:0] x487 ,
input [7:0] x488 ,
input [7:0] x489 ,
input [7:0] x490 ,
input [7:0] x491 ,
input [7:0] x492 ,
input [7:0] x493 ,
input [7:0] x494 ,
input [7:0] x495 ,
input [7:0] x496 ,
input [7:0] x497 ,
input [7:0] x498 ,
input [7:0] x499 ,
input [7:0] x500 ,
input [7:0] x501 ,
input [7:0] x502 ,
input [7:0] x503 ,
input [7:0] x504 ,
input [7:0] x505 ,
input [7:0] x506 ,
input [7:0] x507 ,
input [7:0] x508 ,
input [7:0] x509 ,
input [7:0] x510 ,
input [7:0] x511 ,
input [7:0] x512 ,
input [7:0] x513 ,
input [7:0] x514 ,
input [7:0] x515 ,
input [7:0] x516 ,
input [7:0] x517 ,
input [7:0] x518 ,
input [7:0] x519 ,
input [7:0] x520 ,
input [7:0] x521 ,
input [7:0] x522 ,
input [7:0] x523 ,
input [7:0] x524 ,
input [7:0] x525 ,
input [7:0] x526 ,
input [7:0] x527 ,
input [7:0] x528 ,
input [7:0] x529 ,
input [7:0] x530 ,
input [7:0] x531 ,
input [7:0] x532 ,
input [7:0] x533 ,
input [7:0] x534 ,
input [7:0] x535 ,
input [7:0] x536 ,
input [7:0] x537 ,
input [7:0] x538 ,
input [7:0] x539 ,
input [7:0] x540 ,
input [7:0] x541 ,
input [7:0] x542 ,
input [7:0] x543 ,
input [7:0] x544 ,
input [7:0] x545 ,
input [7:0] x546 ,
input [7:0] x547 ,
input [7:0] x548 ,
input [7:0] x549 ,
input [7:0] x550 ,
input [7:0] x551 ,
input [7:0] x552 ,
input [7:0] x553 ,
input [7:0] x554 ,
input [7:0] x555 ,
input [7:0] x556 ,
input [7:0] x557 ,
input [7:0] x558 ,
input [7:0] x559 ,
input [7:0] x560 ,
input [7:0] x561 ,
input [7:0] x562 ,
input [7:0] x563 ,
input [7:0] x564 ,
input [7:0] x565 ,
input [7:0] x566 ,
input [7:0] x567 ,
input [7:0] x568 ,
input [7:0] x569 ,
input [7:0] x570 ,
input [7:0] x571 ,
input [7:0] x572 ,
input [7:0] x573 ,
input [7:0] x574 ,
input [7:0] x575 ,
input [7:0] x576 ,
input [7:0] x577 ,
input [7:0] x578 ,
input [7:0] x579 ,
input [7:0] x580 ,
input [7:0] x581 ,
input [7:0] x582 ,
input [7:0] x583 ,
input [7:0] x584 ,
input [7:0] x585 ,
input [7:0] x586 ,
input [7:0] x587 ,
input [7:0] x588 ,
input [7:0] x589 ,
input [7:0] x590 ,
input [7:0] x591 ,
input [7:0] x592 ,
input [7:0] x593 ,
input [7:0] x594 ,
input [7:0] x595 ,
input [7:0] x596 ,
input [7:0] x597 ,
input [7:0] x598 ,
input [7:0] x599 ,
input [7:0] x600 ,
input [7:0] x601 ,
input [7:0] x602 ,
input [7:0] x603 ,
input [7:0] x604 ,
input [7:0] x605 ,
input [7:0] x606 ,
input [7:0] x607 ,
input [7:0] x608 ,
input [7:0] x609 ,
input [7:0] x610 ,
input [7:0] x611 ,
input [7:0] x612 ,
input [7:0] x613 ,
input [7:0] x614 ,
input [7:0] x615 ,
input [7:0] x616 ,
input [7:0] x617 ,
input [7:0] x618 ,
input [7:0] x619 ,
input [7:0] x620 ,
input [7:0] x621 ,
input [7:0] x622 ,
input [7:0] x623 ,
input [7:0] x624 ,
input [7:0] x625 ,
input [7:0] x626 ,
input [7:0] x627 ,
input [7:0] x628 ,
input [7:0] x629 ,
input [7:0] x630 ,
input [7:0] x631 ,
input [7:0] x632 ,
input [7:0] x633 ,
input [7:0] x634 ,
input [7:0] x635 ,
input [7:0] x636 ,
input [7:0] x637 ,
input [7:0] x638 ,
input [7:0] x639 ,
input [7:0] x640 ,
input [7:0] x641 ,
input [7:0] x642 ,
input [7:0] x643 ,
input [7:0] x644 ,
input [7:0] x645 ,
input [7:0] x646 ,
input [7:0] x647 ,
input [7:0] x648 ,
input [7:0] x649 ,
input [7:0] x650 ,
input [7:0] x651 ,
input [7:0] x652 ,
input [7:0] x653 ,
input [7:0] x654 ,
input [7:0] x655 ,
input [7:0] x656 ,
input [7:0] x657 ,
input [7:0] x658 ,
input [7:0] x659 ,
input [7:0] x660 ,
input [7:0] x661 ,
input [7:0] x662 ,
input [7:0] x663 ,
input [7:0] x664 ,
input [7:0] x665 ,
input [7:0] x666 ,
input [7:0] x667 ,
input [7:0] x668 ,
input [7:0] x669 ,
input [7:0] x670 ,
input [7:0] x671 ,
input [7:0] x672 ,
input [7:0] x673 ,
input [7:0] x674 ,
input [7:0] x675 ,
input [7:0] x676 ,
input [7:0] x677 ,
input [7:0] x678 ,
input [7:0] x679 ,
input [7:0] x680 ,
input [7:0] x681 ,
input [7:0] x682 ,
input [7:0] x683 ,
input [7:0] x684 ,
input [7:0] x685 ,
input [7:0] x686 ,
input [7:0] x687 ,
input [7:0] x688 ,
input [7:0] x689 ,
input [7:0] x690 ,
input [7:0] x691 ,
input [7:0] x692 ,
input [7:0] x693 ,
input [7:0] x694 ,
input [7:0] x695 ,
input [7:0] x696 ,
input [7:0] x697 ,
input [7:0] x698 ,
input [7:0] x699 ,
input [7:0] x700 ,
input [7:0] x701 ,
input [7:0] x702 ,
input [7:0] x703 ,
input [7:0] x704 ,
input [7:0] x705 ,
input [7:0] x706 ,
input [7:0] x707 ,
input [7:0] x708 ,
input [7:0] x709 ,
input [7:0] x710 ,
input [7:0] x711 ,
input [7:0] x712 ,
input [7:0] x713 ,
input [7:0] x714 ,
input [7:0] x715 ,
input [7:0] x716 ,
input [7:0] x717 ,
input [7:0] x718 ,
input [7:0] x719 ,
input [7:0] x720 ,
input [7:0] x721 ,
input [7:0] x722 ,
input [7:0] x723 ,
input [7:0] x724 ,
input [7:0] x725 ,
input [7:0] x726 ,
input [7:0] x727 ,
input [7:0] x728 ,
input [7:0] x729 ,
input [7:0] x730 ,
input [7:0] x731 ,
input [7:0] x732 ,
input [7:0] x733 ,
input [7:0] x734 ,
input [7:0] x735 ,
input [7:0] x736 ,
input [7:0] x737 ,
input [7:0] x738 ,
input [7:0] x739 ,
input [7:0] x740 ,
input [7:0] x741 ,
input [7:0] x742 ,
input [7:0] x743 ,
input [7:0] x744 ,
input [7:0] x745 ,
input [7:0] x746 ,
input [7:0] x747 ,
input [7:0] x748 ,
input [7:0] x749 ,
input [7:0] x750 ,
input [7:0] x751 ,
input [7:0] x752 ,
input [7:0] x753 ,
input [7:0] x754 ,
input [7:0] x755 ,
input [7:0] x756 ,
input [7:0] x757 ,
input [7:0] x758 ,
input [7:0] x759 ,
input [7:0] x760 ,
input [7:0] x761 ,
input [7:0] x762 ,
input [7:0] x763 ,
input [7:0] x764 ,
input [7:0] x765 ,
input [7:0] x766 ,
input [7:0] x767 ,
input [7:0] x768 ,
input [7:0] x769 ,
input [7:0] x770 ,
input [7:0] x771 ,
input [7:0] x772 ,
input [7:0] x773 ,
input [7:0] x774 ,
input [7:0] x775 ,
input [7:0] x776 ,
input [7:0] x777 ,
input [7:0] x778 ,
input [7:0] x779 ,
input [7:0] x780 ,
input [7:0] x781 ,
input [7:0] x782 ,
input [7:0] x783 ,
input [7:0] x784 ,
input [7:0] x785 ,
input [7:0] x786 ,
input [7:0] x787 ,
input [7:0] x788 ,
input [7:0] x789 ,
input [7:0] x790 ,
input [7:0] x791 ,
input [7:0] x792 ,
input [7:0] x793 ,
input [7:0] x794 ,
input [7:0] x795 ,
input [7:0] x796 ,
input [7:0] x797 ,
input [7:0] x798 ,
input [7:0] x799 ,
input [7:0] x800 ,
input [7:0] x801 ,
input [7:0] x802 ,
input [7:0] x803 ,
input [7:0] x804 ,
input [7:0] x805 ,
input [7:0] x806 ,
input [7:0] x807 ,
input [7:0] x808 ,
input [7:0] x809 ,
input [7:0] x810 ,
input [7:0] x811 ,
input [7:0] x812 ,
input [7:0] x813 ,
input [7:0] x814 ,
input [7:0] x815 ,
input [7:0] x816 ,
input [7:0] x817 ,
input [7:0] x818 ,
input [7:0] x819 ,
input [7:0] x820 ,
input [7:0] x821 ,
input [7:0] x822 ,
input [7:0] x823 ,
input [7:0] x824 ,
input [7:0] x825 ,
input [7:0] x826 ,
input [7:0] x827 ,
input [7:0] x828 ,
input [7:0] x829 ,
input [7:0] x830 ,
input [7:0] x831 ,
input [7:0] x832 ,
input [7:0] x833 ,
input [7:0] x834 ,
input [7:0] x835 ,
input [7:0] x836 ,
input [7:0] x837 ,
input [7:0] x838 ,
input [7:0] x839 ,
input [7:0] x840 ,
input [7:0] x841 ,
input [7:0] x842 ,
input [7:0] x843 ,
input [7:0] x844 ,
input [7:0] x845 ,
input [7:0] x846 ,
input [7:0] x847 ,
input [7:0] x848 ,
input [7:0] x849 ,
input [7:0] x850 ,
input [7:0] x851 ,
input [7:0] x852 ,
input [7:0] x853 ,
input [7:0] x854 ,
input [7:0] x855 ,
input [7:0] x856 ,
input [7:0] x857 ,
input [7:0] x858 ,
input [7:0] x859 ,
input [7:0] x860 ,
input [7:0] x861 ,
input [7:0] x862 ,
input [7:0] x863 ,
input [7:0] x864 ,
input [7:0] x865 ,
input [7:0] x866 ,
input [7:0] x867 ,
input [7:0] x868 ,
input [7:0] x869 ,
input [7:0] x870 ,
input [7:0] x871 ,
input [7:0] x872 ,
input [7:0] x873 ,
input [7:0] x874 ,
input [7:0] x875 ,
input [7:0] x876 ,
input [7:0] x877 ,
input [7:0] x878 ,
input [7:0] x879 ,
input [7:0] x880 ,
input [7:0] x881 ,
input [7:0] x882 ,
input [7:0] x883 ,
input [7:0] x884 ,
input [7:0] x885 ,
input [7:0] x886 ,
input [7:0] x887 ,
input [7:0] x888 ,
input [7:0] x889 ,
input [7:0] x890 ,
input [7:0] x891 ,
input [7:0] x892 ,
input [7:0] x893 ,
input [7:0] x894 ,
input [7:0] x895 ,
input [7:0] x896 ,
input [7:0] x897 ,
input [7:0] x898 ,
input [7:0] x899 ,
input [7:0] x900 ,
input [7:0] x901 ,
input [7:0] x902 ,
input [7:0] x903 ,
input [7:0] x904 ,
input [7:0] x905 ,
input [7:0] x906 ,
input [7:0] x907 ,
input [7:0] x908 ,
input [7:0] x909 ,
input [7:0] x910 ,
input [7:0] x911 ,
input [7:0] x912 ,
input [7:0] x913 ,
input [7:0] x914 ,
input [7:0] x915 ,
input [7:0] x916 ,
input [7:0] x917 ,
input [7:0] x918 ,
input [7:0] x919 ,
input [7:0] x920 ,
input [7:0] x921 ,
input [7:0] x922 ,
input [7:0] x923 ,
input [7:0] x924 ,
input [7:0] x925 ,
input [7:0] x926 ,
input [7:0] x927 ,
input [7:0] x928 ,
input [7:0] x929 ,
input [7:0] x930 ,
input [7:0] x931 ,
input [7:0] x932 ,
input [7:0] x933 ,
input [7:0] x934 ,
input [7:0] x935 ,
input [7:0] x936 ,
input [7:0] x937 ,
input [7:0] x938 ,
input [7:0] x939 ,
input [7:0] x940 ,
input [7:0] x941 ,
input [7:0] x942 ,
input [7:0] x943 ,
input [7:0] x944 ,
input [7:0] x945 ,
input [7:0] x946 ,
input [7:0] x947 ,
input [7:0] x948 ,
input [7:0] x949 ,
input [7:0] x950 ,
input [7:0] x951 ,
input [7:0] x952 ,
input [7:0] x953 ,
input [7:0] x954 ,
input [7:0] x955 ,
input [7:0] x956 ,
input [7:0] x957 ,
input [7:0] x958 ,
input [7:0] x959 ,
input [7:0] x960 ,
input [7:0] x961 ,
input [7:0] x962 ,
input [7:0] x963 ,
input [7:0] x964 ,
input [7:0] x965 ,
input [7:0] x966 ,
input [7:0] x967 ,
input [7:0] x968 ,
input [7:0] x969 ,
input [7:0] x970 ,
input [7:0] x971 ,
input [7:0] x972 ,
input [7:0] x973 ,
input [7:0] x974 ,
input [7:0] x975 ,
input [7:0] x976 ,
input [7:0] x977 ,
input [7:0] x978 ,
input [7:0] x979 ,
input [7:0] x980 ,
input [7:0] x981 ,
input [7:0] x982 ,
input [7:0] x983 ,
input [7:0] x984 ,
input [7:0] x985 ,
input [7:0] x986 ,
input [7:0] x987 ,
input [7:0] x988 ,
input [7:0] x989 ,
input [7:0] x990 ,
input [7:0] x991 ,
input [7:0] x992 ,
input [7:0] x993 ,
input [7:0] x994 ,
input [7:0] x995 ,
input [7:0] x996 ,
input [7:0] x997 ,
input [7:0] x998 ,
input [7:0] x999 ,
input [7:0] x1000 ,
input [7:0] x1001 ,
input [7:0] x1002 ,
input [7:0] x1003 ,
input [7:0] x1004 ,
input [7:0] x1005 ,
input [7:0] x1006 ,
input [7:0] x1007 ,
input [7:0] x1008 ,
input [7:0] x1009 ,
input [7:0] x1010 ,
input [7:0] x1011 ,
input [7:0] x1012 ,
input [7:0] x1013 ,
input [7:0] x1014 ,
input [7:0] x1015 ,
input [7:0] x1016 ,
input [7:0] x1017 ,
input [7:0] x1018 ,
input [7:0] x1019 ,
input [7:0] x1020 ,
input [7:0] x1021 ,
input [7:0] x1022 ,
input [7:0] x1023 ,
input [7:0] x1024 ,
input [7:0] x1025 ,
input [7:0] x1026 ,
input [7:0] x1027 ,
input [7:0] x1028 ,
input [7:0] x1029 ,
input [7:0] x1030 ,
input [7:0] x1031 ,
input [7:0] x1032 ,
input [7:0] x1033 ,
input [7:0] x1034 ,
input [7:0] x1035 ,
input [7:0] x1036 ,
input [7:0] x1037 ,
input [7:0] x1038 ,
input [7:0] x1039 ,
input [7:0] x1040 ,
input [7:0] x1041 ,
input [7:0] x1042 ,
input [7:0] x1043 ,
input [7:0] x1044 ,
input [7:0] x1045 ,
input [7:0] x1046 ,
input [7:0] x1047 ,
input [7:0] x1048 ,
input [7:0] x1049 ,
input [7:0] x1050 ,
input [7:0] x1051 ,
input [7:0] x1052 ,
input [7:0] x1053 ,
input [7:0] x1054 ,
input [7:0] x1055 ,
input [7:0] x1056 ,
input [7:0] x1057 ,
input [7:0] x1058 ,
input [7:0] x1059 ,
input [7:0] x1060 ,
input [7:0] x1061 ,
input [7:0] x1062 ,
input [7:0] x1063 ,
input [7:0] x1064 ,
input [7:0] x1065 ,
input [7:0] x1066 ,
input [7:0] x1067 ,
input [7:0] x1068 ,
input [7:0] x1069 ,
input [7:0] x1070 ,
input [7:0] x1071 ,
input [7:0] x1072 ,
input [7:0] x1073 ,
input [7:0] x1074 ,
input [7:0] x1075 ,
input [7:0] x1076 ,
input [7:0] x1077 ,
input [7:0] x1078 ,
input [7:0] x1079 ,
input [7:0] x1080 ,
input [7:0] x1081 ,
input [7:0] x1082 ,
input [7:0] x1083 ,
input [7:0] x1084 ,
input [7:0] x1085 ,
input [7:0] x1086 ,
input [7:0] x1087 ,
input [7:0] x1088 ,
input [7:0] x1089 ,
input [7:0] x1090 ,
input [7:0] x1091 ,
input [7:0] x1092 ,
input [7:0] x1093 ,
input [7:0] x1094 ,
input [7:0] x1095 ,
input [7:0] x1096 ,
input [7:0] x1097 ,
input [7:0] x1098 ,
input [7:0] x1099 ,
input [7:0] x1100 ,
input [7:0] x1101 ,
input [7:0] x1102 ,
input [7:0] x1103 ,
input [7:0] x1104 ,
input [7:0] x1105 ,
input [7:0] x1106 ,
input [7:0] x1107 ,
input [7:0] x1108 ,
input [7:0] x1109 ,
input [7:0] x1110 ,
input [7:0] x1111 ,
input [7:0] x1112 ,
input [7:0] x1113 ,
input [7:0] x1114 ,
input [7:0] x1115 ,
input [7:0] x1116 ,
input [7:0] x1117 ,
input [7:0] x1118 ,
input [7:0] x1119 ,
input [7:0] x1120 ,
input [7:0] x1121 ,
input [7:0] x1122 ,
input [7:0] x1123 ,
input [7:0] x1124 ,
input [7:0] x1125 ,
input [7:0] x1126 ,
input [7:0] x1127 ,
input [7:0] x1128 ,
input [7:0] x1129 ,
input [7:0] x1130 ,
input [7:0] x1131 ,
input [7:0] x1132 ,
input [7:0] x1133 ,
input [7:0] x1134 ,
input [7:0] x1135 ,
input [7:0] x1136 ,
input [7:0] x1137 ,
input [7:0] x1138 ,
input [7:0] x1139 ,
input [7:0] x1140 ,
input [7:0] x1141 ,
input [7:0] x1142 ,
input [7:0] x1143 ,
input [7:0] x1144 ,
input [7:0] x1145 ,
input [7:0] x1146 ,
input [7:0] x1147 ,
input [7:0] x1148 ,
input [7:0] x1149 ,
input [7:0] x1150 ,
input [7:0] x1151 ,
input [7:0] x1152 ,
input [7:0] x1153 ,
input [7:0] x1154 ,
input [7:0] x1155 ,
input [7:0] x1156 ,
input [7:0] x1157 ,
input [7:0] x1158 ,
input [7:0] x1159 ,
input [7:0] x1160 ,
input [7:0] x1161 ,
input [7:0] x1162 ,
input [7:0] x1163 ,
input [7:0] x1164 ,
input [7:0] x1165 ,
input [7:0] x1166 ,
input [7:0] x1167 ,
input [7:0] x1168 ,
input [7:0] x1169 ,
input [7:0] x1170 ,
input [7:0] x1171 ,
input [7:0] x1172 ,
input [7:0] x1173 ,
input [7:0] x1174 ,
input [7:0] x1175 ,
input [7:0] x1176 ,
input [7:0] x1177 ,
input [7:0] x1178 ,
input [7:0] x1179 ,
input [7:0] x1180 ,
input [7:0] x1181 ,
input [7:0] x1182 ,
input [7:0] x1183 ,
input [7:0] x1184 ,
input [7:0] x1185 ,
input [7:0] x1186 ,
input [7:0] x1187 ,
input [7:0] x1188 ,
input [7:0] x1189 ,
input [7:0] x1190 ,
input [7:0] x1191 ,
input [7:0] x1192 ,
input [7:0] x1193 ,
input [7:0] x1194 ,
input [7:0] x1195 ,
input [7:0] x1196 ,
input [7:0] x1197 ,
input [7:0] x1198 ,
input [7:0] x1199 ,
input [7:0] x1200 ,
input [7:0] x1201 ,
input [7:0] x1202 ,
input [7:0] x1203 ,
input [7:0] x1204 ,
input [7:0] x1205 ,
input [7:0] x1206 ,
input [7:0] x1207 ,
input [7:0] x1208 ,
input [7:0] x1209 ,
input [7:0] x1210 ,
input [7:0] x1211 ,
input [7:0] x1212 ,
input [7:0] x1213 ,
input [7:0] x1214 ,
input [7:0] x1215 ,
input [7:0] x1216 ,
input [7:0] x1217 ,
input [7:0] x1218 ,
input [7:0] x1219 ,
input [7:0] x1220 ,
input [7:0] x1221 ,
input [7:0] x1222 ,
input [7:0] x1223 ,
input [7:0] x1224 ,
input [7:0] x1225 ,
input [7:0] x1226 ,
input [7:0] x1227 ,
input [7:0] x1228 ,
input [7:0] x1229 ,
input [7:0] x1230 ,
input [7:0] x1231 ,
input [7:0] x1232 ,
input [7:0] x1233 ,
input [7:0] x1234 ,
input [7:0] x1235 ,
input [7:0] x1236 ,
input [7:0] x1237 ,
input [7:0] x1238 ,
input [7:0] x1239 ,
input [7:0] x1240 ,
input [7:0] x1241 ,
input [7:0] x1242 ,
input [7:0] x1243 ,
input [7:0] x1244 ,
input [7:0] x1245 ,
input [7:0] x1246 ,
input [7:0] x1247 ,
input [7:0] x1248 ,
input [7:0] x1249 ,
input [7:0] x1250 ,
input [7:0] x1251 ,
input [7:0] x1252 ,
input [7:0] x1253 ,
input [7:0] x1254 ,
input [7:0] x1255 ,
input [7:0] x1256 ,
input [7:0] x1257 ,
input [7:0] x1258 ,
input [7:0] x1259 ,
input [7:0] x1260 ,
input [7:0] x1261 ,
input [7:0] x1262 ,
input [7:0] x1263 ,
input [7:0] x1264 ,
input [7:0] x1265 ,
input [7:0] x1266 ,
input [7:0] x1267 ,
input [7:0] x1268 ,
input [7:0] x1269 ,
input [7:0] x1270 ,
input [7:0] x1271 ,
input [7:0] x1272 ,
input [7:0] x1273 ,
input [7:0] x1274 ,
input [7:0] x1275 ,
input [7:0] x1276 ,
input [7:0] x1277 ,
input [7:0] x1278 ,
input [7:0] x1279 ,
input [7:0] x1280 ,
input [7:0] x1281 ,
input [7:0] x1282 ,
input [7:0] x1283 ,
input [7:0] x1284 ,
input [7:0] x1285 ,
input [7:0] x1286 ,
input [7:0] x1287 ,
input [7:0] x1288 ,
input [7:0] x1289 ,
input [7:0] x1290 ,
input [7:0] x1291 ,
input [7:0] x1292 ,
input [7:0] x1293 ,
input [7:0] x1294 ,
input [7:0] x1295 ,
input [7:0] x1296 ,
input [7:0] x1297 ,
input [7:0] x1298 ,
input [7:0] x1299 ,
input [7:0] x1300 ,
input [7:0] x1301 ,
input [7:0] x1302 ,
input [7:0] x1303 ,
input [7:0] x1304 ,
input [7:0] x1305 ,
input [7:0] x1306 ,
input [7:0] x1307 ,
input [7:0] x1308 ,
input [7:0] x1309 ,
input [7:0] x1310 ,
input [7:0] x1311 ,
input [7:0] x1312 ,
input [7:0] x1313 ,
input [7:0] x1314 ,
input [7:0] x1315 ,
input [7:0] x1316 ,
input [7:0] x1317 ,
input [7:0] x1318 ,
input [7:0] x1319 ,
input [7:0] x1320 ,
input [7:0] x1321 ,
input [7:0] x1322 ,
input [7:0] x1323 ,
input [7:0] x1324 ,
input [7:0] x1325 ,
input [7:0] x1326 ,
input [7:0] x1327 ,
input [7:0] x1328 ,
input [7:0] x1329 ,
input [7:0] x1330 ,
input [7:0] x1331 ,
input [7:0] x1332 ,
input [7:0] x1333 ,
input [7:0] x1334 ,
input [7:0] x1335 ,
input [7:0] x1336 ,
input [7:0] x1337 ,
input [7:0] x1338 ,
input [7:0] x1339 ,
input [7:0] x1340 ,
input [7:0] x1341 ,
input [7:0] x1342 ,
input [7:0] x1343 ,
input [7:0] x1344 ,
input [7:0] x1345 ,
input [7:0] x1346 ,
input [7:0] x1347 ,
input [7:0] x1348 ,
input [7:0] x1349 ,
input [7:0] x1350 ,
input [7:0] x1351 ,
input [7:0] x1352 ,
input [7:0] x1353 ,
input [7:0] x1354 ,
input [7:0] x1355 ,
input [7:0] x1356 ,
input [7:0] x1357 ,
input [7:0] x1358 ,
input [7:0] x1359 ,
input [7:0] x1360 ,
input [7:0] x1361 ,
input [7:0] x1362 ,
input [7:0] x1363 ,
input [7:0] x1364 ,
input [7:0] x1365 ,
input [7:0] x1366 ,
input [7:0] x1367 ,
input [7:0] x1368 ,
input [7:0] x1369 ,
input [7:0] x1370 ,
input [7:0] x1371 ,
input [7:0] x1372 ,
input [7:0] x1373 ,
input [7:0] x1374 ,
input [7:0] x1375 ,
input [7:0] x1376 ,
input [7:0] x1377 ,
input [7:0] x1378 ,
input [7:0] x1379 ,
input [7:0] x1380 ,
input [7:0] x1381 ,
input [7:0] x1382 ,
input [7:0] x1383 ,
input [7:0] x1384 ,
input [7:0] x1385 ,
input [7:0] x1386 ,
input [7:0] x1387 ,
input [7:0] x1388 ,
input [7:0] x1389 ,
input [7:0] x1390 ,
input [7:0] x1391 ,
input [7:0] x1392 ,
input [7:0] x1393 ,
input [7:0] x1394 ,
input [7:0] x1395 ,
input [7:0] x1396 ,
input [7:0] x1397 ,
input [7:0] x1398 ,
input [7:0] x1399 ,
input [7:0] x1400 ,
input [7:0] x1401 ,
input [7:0] x1402 ,
input [7:0] x1403 ,
input [7:0] x1404 ,
input [7:0] x1405 ,
input [7:0] x1406 ,
input [7:0] x1407 ,
input [7:0] x1408 ,
input [7:0] x1409 ,
input [7:0] x1410 ,
input [7:0] x1411 ,
input [7:0] x1412 ,
input [7:0] x1413 ,
input [7:0] x1414 ,
input [7:0] x1415 ,
input [7:0] x1416 ,
input [7:0] x1417 ,
input [7:0] x1418 ,
input [7:0] x1419 ,
input [7:0] x1420 ,
input [7:0] x1421 ,
input [7:0] x1422 ,
input [7:0] x1423 ,
input [7:0] x1424 ,
input [7:0] x1425 ,
input [7:0] x1426 ,
input [7:0] x1427 ,
input [7:0] x1428 ,
input [7:0] x1429 ,
input [7:0] x1430 ,
input [7:0] x1431 ,
input [7:0] x1432 ,
input [7:0] x1433 ,
input [7:0] x1434 ,
input [7:0] x1435 ,
input [7:0] x1436 ,
input [7:0] x1437 ,
input [7:0] x1438 ,
input [7:0] x1439 ,
input [7:0] x1440 ,
input [7:0] x1441 ,
input [7:0] x1442 ,
input [7:0] x1443 ,
input [7:0] x1444 ,
input [7:0] x1445 ,
input [7:0] x1446 ,
input [7:0] x1447 ,
input [7:0] x1448 ,
input [7:0] x1449 ,
input [7:0] x1450 ,
input [7:0] x1451 ,
input [7:0] x1452 ,
input [7:0] x1453 ,
input [7:0] x1454 ,
input [7:0] x1455 ,
input [7:0] x1456 ,
input [7:0] x1457 ,
input [7:0] x1458 ,
input [7:0] x1459 ,
input [7:0] x1460 ,
input [7:0] x1461 ,
input [7:0] x1462 ,
input [7:0] x1463 ,
input [7:0] x1464 ,
input [7:0] x1465 ,
input [7:0] x1466 ,
input [7:0] x1467 ,
input [7:0] x1468 ,
input [7:0] x1469 ,
input [7:0] x1470 ,
input [7:0] x1471 ,
input [7:0] x1472 ,
input [7:0] x1473 ,
input [7:0] x1474 ,
input [7:0] x1475 ,
input [7:0] x1476 ,
input [7:0] x1477 ,
input [7:0] x1478 ,
input [7:0] x1479 ,
input [7:0] x1480 ,
input [7:0] x1481 ,
input [7:0] x1482 ,
input [7:0] x1483 ,
input [7:0] x1484 ,
input [7:0] x1485 ,
input [7:0] x1486 ,
input [7:0] x1487 ,
input [7:0] x1488 ,
input [7:0] x1489 ,
input [7:0] x1490 ,
input [7:0] x1491 ,
input [7:0] x1492 ,
input [7:0] x1493 ,
input [7:0] x1494 ,
input [7:0] x1495 ,
input [7:0] x1496 ,
input [7:0] x1497 ,
input [7:0] x1498 ,
input [7:0] x1499 ,
input [7:0] x1500 ,
input [7:0] x1501 ,
input [7:0] x1502 ,
input [7:0] x1503 ,
input [7:0] x1504 ,
input [7:0] x1505 ,
input [7:0] x1506 ,
input [7:0] x1507 ,
input [7:0] x1508 ,
input [7:0] x1509 ,
input [7:0] x1510 ,
input [7:0] x1511 ,
input [7:0] x1512 ,
input [7:0] x1513 ,
input [7:0] x1514 ,
input [7:0] x1515 ,
input [7:0] x1516 ,
input [7:0] x1517 ,
input [7:0] x1518 ,
input [7:0] x1519 ,
input [7:0] x1520 ,
input [7:0] x1521 ,
input [7:0] x1522 ,
input [7:0] x1523 ,
input [7:0] x1524 ,
input [7:0] x1525 ,
input [7:0] x1526 ,
input [7:0] x1527 ,
input [7:0] x1528 ,
input [7:0] x1529 ,
input [7:0] x1530 ,
input [7:0] x1531 ,
input [7:0] x1532 ,
input [7:0] x1533 ,
input [7:0] x1534 ,
input [7:0] x1535 ,
input [7:0] x1536 ,
input [7:0] x1537 ,
input [7:0] x1538 ,
input [7:0] x1539 ,
input [7:0] x1540 ,
input [7:0] x1541 ,
input [7:0] x1542 ,
input [7:0] x1543 ,
input [7:0] x1544 ,
input [7:0] x1545 ,
input [7:0] x1546 ,
input [7:0] x1547 ,
input [7:0] x1548 ,
input [7:0] x1549 ,
input [7:0] x1550 ,
input [7:0] x1551 ,
input [7:0] x1552 ,
input [7:0] x1553 ,
input [7:0] x1554 ,
input [7:0] x1555 ,
input [7:0] x1556 ,
input [7:0] x1557 ,
input [7:0] x1558 ,
input [7:0] x1559 ,
input [7:0] x1560 ,
input [7:0] x1561 ,
input [7:0] x1562 ,
input [7:0] x1563 ,
input [7:0] x1564 ,
input [7:0] x1565 ,
input [7:0] x1566 ,
input [7:0] x1567 ,
input [7:0] x1568 ,
input [7:0] x1569 ,
input [7:0] x1570 ,
input [7:0] x1571 ,
input [7:0] x1572 ,
input [7:0] x1573 ,
input [7:0] x1574 ,
input [7:0] x1575 ,
input [7:0] x1576 ,
input [7:0] x1577 ,
input [7:0] x1578 ,
input [7:0] x1579 ,
input [7:0] x1580 ,
input [7:0] x1581 ,
input [7:0] x1582 ,
input [7:0] x1583 ,
input [7:0] x1584 ,
input [7:0] x1585 ,
input [7:0] x1586 ,
input [7:0] x1587 ,
input [7:0] x1588 ,
input [7:0] x1589 ,
input [7:0] x1590 ,
input [7:0] x1591 ,
input [7:0] x1592 ,
input [7:0] x1593 ,
input [7:0] x1594 ,
input [7:0] x1595 ,
input [7:0] x1596 ,
input [7:0] x1597 ,
input [7:0] x1598 ,
input [7:0] x1599 ,
input [7:0] x1600 ,
input [7:0] x1601 ,
input [7:0] x1602 ,
input [7:0] x1603 ,
input [7:0] x1604 ,
input [7:0] x1605 ,
input [7:0] x1606 ,
input [7:0] x1607 ,
input [7:0] x1608 ,
input [7:0] x1609 ,
input [7:0] x1610 ,
input [7:0] x1611 ,
input [7:0] x1612 ,
input [7:0] x1613 ,
input [7:0] x1614 ,
input [7:0] x1615 ,
input [7:0] x1616 ,
input [7:0] x1617 ,
input [7:0] x1618 ,
input [7:0] x1619 ,
input [7:0] x1620 ,
input [7:0] x1621 ,
input [7:0] x1622 ,
input [7:0] x1623 ,
input [7:0] x1624 ,
input [7:0] x1625 ,
input [7:0] x1626 ,
input [7:0] x1627 ,
input [7:0] x1628 ,
input [7:0] x1629 ,
input [7:0] x1630 ,
input [7:0] x1631 ,
input [7:0] x1632 ,
input [7:0] x1633 ,
input [7:0] x1634 ,
input [7:0] x1635 ,
input [7:0] x1636 ,
input [7:0] x1637 ,
input [7:0] x1638 ,
input [7:0] x1639 ,
input [7:0] x1640 ,
input [7:0] x1641 ,
input [7:0] x1642 ,
input [7:0] x1643 ,
input [7:0] x1644 ,
input [7:0] x1645 ,
input [7:0] x1646 ,
input [7:0] x1647 ,
input [7:0] x1648 ,
input [7:0] x1649 ,
input [7:0] x1650 ,
input [7:0] x1651 ,
input [7:0] x1652 ,
input [7:0] x1653 ,
input [7:0] x1654 ,
input [7:0] x1655 ,
input [7:0] x1656 ,
input [7:0] x1657 ,
input [7:0] x1658 ,
input [7:0] x1659 ,
input [7:0] x1660 ,
input [7:0] x1661 ,
input [7:0] x1662 ,
input [7:0] x1663 ,
input [7:0] x1664 ,
input [7:0] x1665 ,
input [7:0] x1666 ,
input [7:0] x1667 ,
input [7:0] x1668 ,
input [7:0] x1669 ,
input [7:0] x1670 ,
input [7:0] x1671 ,
input [7:0] x1672 ,
input [7:0] x1673 ,
input [7:0] x1674 ,
input [7:0] x1675 ,
input [7:0] x1676 ,
input [7:0] x1677 ,
input [7:0] x1678 ,
input [7:0] x1679 ,
input [7:0] x1680 ,
input [7:0] x1681 ,
input [7:0] x1682 ,
input [7:0] x1683 ,
input [7:0] x1684 ,
input [7:0] x1685 ,
input [7:0] x1686 ,
input [7:0] x1687 ,
input [7:0] x1688 ,
input [7:0] x1689 ,
input [7:0] x1690 ,
input [7:0] x1691 ,
input [7:0] x1692 ,
input [7:0] x1693 ,
input [7:0] x1694 ,
input [7:0] x1695 ,
input [7:0] x1696 ,
input [7:0] x1697 ,
input [7:0] x1698 ,
input [7:0] x1699 ,
input [7:0] x1700 ,
input [7:0] x1701 ,
input [7:0] x1702 ,
input [7:0] x1703 ,
input [7:0] x1704 ,
input [7:0] x1705 ,
input [7:0] x1706 ,
input [7:0] x1707 ,
input [7:0] x1708 ,
input [7:0] x1709 ,
input [7:0] x1710 ,
input [7:0] x1711 ,
input [7:0] x1712 ,
input [7:0] x1713 ,
input [7:0] x1714 ,
input [7:0] x1715 ,
input [7:0] x1716 ,
input [7:0] x1717 ,
input [7:0] x1718 ,
input [7:0] x1719 ,
input [7:0] x1720 ,
input [7:0] x1721 ,
input [7:0] x1722 ,
input [7:0] x1723 ,
input [7:0] x1724 ,
input [7:0] x1725 ,
input [7:0] x1726 ,
input [7:0] x1727 ,
input [7:0] x1728 ,
input [7:0] x1729 ,
input [7:0] x1730 ,
input [7:0] x1731 ,
input [7:0] x1732 ,
input [7:0] x1733 ,
input [7:0] x1734 ,
input [7:0] x1735 ,
input [7:0] x1736 ,
input [7:0] x1737 ,
input [7:0] x1738 ,
input [7:0] x1739 ,
input [7:0] x1740 ,
input [7:0] x1741 ,
input [7:0] x1742 ,
input [7:0] x1743 ,
input [7:0] x1744 ,
input [7:0] x1745 ,
input [7:0] x1746 ,
input [7:0] x1747 ,
input [7:0] x1748 ,
input [7:0] x1749 ,
input [7:0] x1750 ,
input [7:0] x1751 ,
input [7:0] x1752 ,
input [7:0] x1753 ,
input [7:0] x1754 ,
input [7:0] x1755 ,
input [7:0] x1756 ,
input [7:0] x1757 ,
input [7:0] x1758 ,
input [7:0] x1759 ,
input [7:0] x1760 ,
input [7:0] x1761 ,
input [7:0] x1762 ,
input [7:0] x1763 ,
input [7:0] x1764 ,
input [7:0] x1765 ,
input [7:0] x1766 ,
input [7:0] x1767 ,
input [7:0] x1768 ,
input [7:0] x1769 ,
input [7:0] x1770 ,
input [7:0] x1771 ,
input [7:0] x1772 ,
input [7:0] x1773 ,
input [7:0] x1774 ,
input [7:0] x1775 ,
input [7:0] x1776 ,
input [7:0] x1777 ,
input [7:0] x1778 ,
input [7:0] x1779 ,
input [7:0] x1780 ,
input [7:0] x1781 ,
input [7:0] x1782 ,
input [7:0] x1783 ,
input [7:0] x1784 ,
input [7:0] x1785 ,
input [7:0] x1786 ,
input [7:0] x1787 ,
input [7:0] x1788 ,
input [7:0] x1789 ,
input [7:0] x1790 ,
input [7:0] x1791 ,
input [7:0] x1792 ,
input [7:0] x1793 ,
input [7:0] x1794 ,
input [7:0] x1795 ,
input [7:0] x1796 ,
input [7:0] x1797 ,
input [7:0] x1798 ,
input [7:0] x1799 ,
input [7:0] x1800 ,
input [7:0] x1801 ,
input [7:0] x1802 ,
input [7:0] x1803 ,
input [7:0] x1804 ,
input [7:0] x1805 ,
input [7:0] x1806 ,
input [7:0] x1807 ,
input [7:0] x1808 ,
input [7:0] x1809 ,
input [7:0] x1810 ,
input [7:0] x1811 ,
input [7:0] x1812 ,
input [7:0] x1813 ,
input [7:0] x1814 ,
input [7:0] x1815 ,
input [7:0] x1816 ,
input [7:0] x1817 ,
input [7:0] x1818 ,
input [7:0] x1819 ,
input [7:0] x1820 ,
input [7:0] x1821 ,
input [7:0] x1822 ,
input [7:0] x1823 ,
input [7:0] x1824 ,
input [7:0] x1825 ,
input [7:0] x1826 ,
input [7:0] x1827 ,
input [7:0] x1828 ,
input [7:0] x1829 ,
input [7:0] x1830 ,
input [7:0] x1831 ,
input [7:0] x1832 ,
input [7:0] x1833 ,
input [7:0] x1834 ,
input [7:0] x1835 ,
input [7:0] x1836 ,
input [7:0] x1837 ,
input [7:0] x1838 ,
input [7:0] x1839 ,
input [7:0] x1840 ,
input [7:0] x1841 ,
input [7:0] x1842 ,
input [7:0] x1843 ,
input [7:0] x1844 ,
input [7:0] x1845 ,
input [7:0] x1846 ,
input [7:0] x1847 ,
input [7:0] x1848 ,
input [7:0] x1849 ,
input [7:0] x1850 ,
input [7:0] x1851 ,
input [7:0] x1852 ,
input [7:0] x1853 ,
input [7:0] x1854 ,
input [7:0] x1855 ,
input [7:0] x1856 ,
input [7:0] x1857 ,
input [7:0] x1858 ,
input [7:0] x1859 ,
input [7:0] x1860 ,
input [7:0] x1861 ,
input [7:0] x1862 ,
input [7:0] x1863 ,
input [7:0] x1864 ,
input [7:0] x1865 ,
input [7:0] x1866 ,
input [7:0] x1867 ,
input [7:0] x1868 ,
input [7:0] x1869 ,
input [7:0] x1870 ,
input [7:0] x1871 ,
input [7:0] x1872 ,
input [7:0] x1873 ,
input [7:0] x1874 ,
input [7:0] x1875 ,
input [7:0] x1876 ,
input [7:0] x1877 ,
input [7:0] x1878 ,
input [7:0] x1879 ,
input [7:0] x1880 ,
input [7:0] x1881 ,
input [7:0] x1882 ,
input [7:0] x1883 ,
input [7:0] x1884 ,
input [7:0] x1885 ,
input [7:0] x1886 ,
input [7:0] x1887 ,
input [7:0] x1888 ,
input [7:0] x1889 ,
input [7:0] x1890 ,
input [7:0] x1891 ,
input [7:0] x1892 ,
input [7:0] x1893 ,
input [7:0] x1894 ,
input [7:0] x1895 ,
input [7:0] x1896 ,
input [7:0] x1897 ,
input [7:0] x1898 ,
input [7:0] x1899 ,
input [7:0] x1900 ,
input [7:0] x1901 ,
input [7:0] x1902 ,
input [7:0] x1903 ,
input [7:0] x1904 ,
input [7:0] x1905 ,
input [7:0] x1906 ,
input [7:0] x1907 ,
input [7:0] x1908 ,
input [7:0] x1909 ,
input [7:0] x1910 ,
input [7:0] x1911 ,
input [7:0] x1912 ,
input [7:0] x1913 ,
input [7:0] x1914 ,
input [7:0] x1915 ,
input [7:0] x1916 ,
input [7:0] x1917 ,
input [7:0] x1918 ,
input [7:0] x1919 ,
input [7:0] x1920 ,
input [7:0] x1921 ,
input [7:0] x1922 ,
input [7:0] x1923 ,
input [7:0] x1924 ,
input [7:0] x1925 ,
input [7:0] x1926 ,
input [7:0] x1927 ,
input [7:0] x1928 ,
input [7:0] x1929 ,
input [7:0] x1930 ,
input [7:0] x1931 ,
input [7:0] x1932 ,
input [7:0] x1933 ,
input [7:0] x1934 ,
input [7:0] x1935 ,
input [7:0] x1936 ,
input [7:0] x1937 ,
input [7:0] x1938 ,
input [7:0] x1939 ,
input [7:0] x1940 ,
input [7:0] x1941 ,
input [7:0] x1942 ,
input [7:0] x1943 ,
input [7:0] x1944 ,
input [7:0] x1945 ,
input [7:0] x1946 ,
input [7:0] x1947 ,
input [7:0] x1948 ,
input [7:0] x1949 ,
input [7:0] x1950 ,
input [7:0] x1951 ,
input [7:0] x1952 ,
input [7:0] x1953 ,
input [7:0] x1954 ,
input [7:0] x1955 ,
input [7:0] x1956 ,
input [7:0] x1957 ,
input [7:0] x1958 ,
input [7:0] x1959 ,
input [7:0] x1960 ,
input [7:0] x1961 ,
input [7:0] x1962 ,
input [7:0] x1963 ,
input [7:0] x1964 ,
input [7:0] x1965 ,
input [7:0] x1966 ,
input [7:0] x1967 ,
input [7:0] x1968 ,
input [7:0] x1969 ,
input [7:0] x1970 ,
input [7:0] x1971 ,
input [7:0] x1972 ,
input [7:0] x1973 ,
input [7:0] x1974 ,
input [7:0] x1975 ,
input [7:0] x1976 ,
input [7:0] x1977 ,
input [7:0] x1978 ,
input [7:0] x1979 ,
input [7:0] x1980 ,
input [7:0] x1981 ,
input [7:0] x1982 ,
input [7:0] x1983 ,
input [7:0] x1984 ,
input [7:0] x1985 ,
input [7:0] x1986 ,
input [7:0] x1987 ,
input [7:0] x1988 ,
input [7:0] x1989 ,
input [7:0] x1990 ,
input [7:0] x1991 ,
input [7:0] x1992 ,
input [7:0] x1993 ,
input [7:0] x1994 ,
input [7:0] x1995 ,
input [7:0] x1996 ,
input [7:0] x1997 ,
input [7:0] x1998 ,
input [7:0] x1999 ,
input [7:0] x2000 ,
input [7:0] x2001 ,
input [7:0] x2002 ,
input [7:0] x2003 ,
input [7:0] x2004 ,
input [7:0] x2005 ,
input [7:0] x2006 ,
input [7:0] x2007 ,
input [7:0] x2008 ,
input [7:0] x2009 ,
input [7:0] x2010 ,
input [7:0] x2011 ,
input [7:0] x2012 ,
input [7:0] x2013 ,
input [7:0] x2014 ,
input [7:0] x2015 ,
input [7:0] x2016 ,
input [7:0] x2017 ,
input [7:0] x2018 ,
input [7:0] x2019 ,
input [7:0] x2020 ,
input [7:0] x2021 ,
input [7:0] x2022 ,
input [7:0] x2023 ,
input [7:0] x2024 ,
input [7:0] x2025 ,
input [7:0] x2026 ,
input [7:0] x2027 ,
input [7:0] x2028 ,
input [7:0] x2029 ,
input [7:0] x2030 ,
input [7:0] x2031 ,
input [7:0] x2032 ,
input [7:0] x2033 ,
input [7:0] x2034 ,
input [7:0] x2035 ,
input [7:0] x2036 ,
input [7:0] x2037 ,
input [7:0] x2038 ,
input [7:0] x2039 ,
input [7:0] x2040 ,
input [7:0] x2041 ,
input [7:0] x2042 ,
input [7:0] x2043 ,
input [7:0] x2044 ,
input [7:0] x2045 ,
input [7:0] x2046 ,
input [7:0] x2047 ,
input [7:0] x2048 ,
input [7:0] x2049 ,
input [7:0] x2050 ,
input [7:0] x2051 ,
input [7:0] x2052 ,
input [7:0] x2053 ,
input [7:0] x2054 ,
input [7:0] x2055 ,
input [7:0] x2056 ,
input [7:0] x2057 ,
input [7:0] x2058 ,
input [7:0] x2059 ,
input [7:0] x2060 ,
input [7:0] x2061 ,
input [7:0] x2062 ,
input [7:0] x2063 ,
input [7:0] x2064 ,
input [7:0] x2065 ,
input [7:0] x2066 ,
input [7:0] x2067 ,
input [7:0] x2068 ,
input [7:0] x2069 ,
input [7:0] x2070 ,
input [7:0] x2071 ,
input [7:0] x2072 ,
input [7:0] x2073 ,
input [7:0] x2074 ,
input [7:0] x2075 ,
input [7:0] x2076 ,
input [7:0] x2077 ,
input [7:0] x2078 ,
input [7:0] x2079 ,
input [7:0] x2080 ,
input [7:0] x2081 ,
input [7:0] x2082 ,
input [7:0] x2083 ,
input [7:0] x2084 ,
input [7:0] x2085 ,
input [7:0] x2086 ,
input [7:0] x2087 ,
input [7:0] x2088 ,
input [7:0] x2089 ,
input [7:0] x2090 ,
input [7:0] x2091 ,
input [7:0] x2092 ,
input [7:0] x2093 ,
input [7:0] x2094 ,
input [7:0] x2095 ,
input [7:0] x2096 ,
input [7:0] x2097 ,
input [7:0] x2098 ,
input [7:0] x2099 ,
input [7:0] x2100 ,
input [7:0] x2101 ,
input [7:0] x2102 ,
input [7:0] x2103 ,
input [7:0] x2104 ,
input [7:0] x2105 ,
input [7:0] x2106 ,
input [7:0] x2107 ,
input [7:0] x2108 ,
input [7:0] x2109 ,
input [7:0] x2110 ,
input [7:0] x2111 ,
input [7:0] x2112 ,
input [7:0] x2113 ,
input [7:0] x2114 ,
input [7:0] x2115 ,
input [7:0] x2116 ,
input [7:0] x2117 ,
input [7:0] x2118 ,
input [7:0] x2119 ,
input [7:0] x2120 ,
input [7:0] x2121 ,
input [7:0] x2122 ,
input [7:0] x2123 ,
input [7:0] x2124 ,
input [7:0] x2125 ,
input [7:0] x2126 ,
input [7:0] x2127 ,
input [7:0] x2128 ,
input [7:0] x2129 ,
input [7:0] x2130 ,
input [7:0] x2131 ,
input [7:0] x2132 ,
input [7:0] x2133 ,
input [7:0] x2134 ,
input [7:0] x2135 ,
input [7:0] x2136 ,
input [7:0] x2137 ,
input [7:0] x2138 ,
input [7:0] x2139 ,
input [7:0] x2140 ,
input [7:0] x2141 ,
input [7:0] x2142 ,
input [7:0] x2143 ,
input [7:0] x2144 ,
input [7:0] x2145 ,
input [7:0] x2146 ,
input [7:0] x2147 ,
input [7:0] x2148 ,
input [7:0] x2149 ,
input [7:0] x2150 ,
input [7:0] x2151 ,
input [7:0] x2152 ,
input [7:0] x2153 ,
input [7:0] x2154 ,
input [7:0] x2155 ,
input [7:0] x2156 ,
input [7:0] x2157 ,
input [7:0] x2158 ,
input [7:0] x2159 ,
input [7:0] x2160 ,
input [7:0] x2161 ,
input [7:0] x2162 ,
input [7:0] x2163 ,
input [7:0] x2164 ,
input [7:0] x2165 ,
input [7:0] x2166 ,
input [7:0] x2167 ,
input [7:0] x2168 ,
input [7:0] x2169 ,
input [7:0] x2170 ,
input [7:0] x2171 ,
input [7:0] x2172 ,
input [7:0] x2173 ,
input [7:0] x2174 ,
input [7:0] x2175 ,
input [7:0] x2176 ,
input [7:0] x2177 ,
input [7:0] x2178 ,
input [7:0] x2179 ,
input [7:0] x2180 ,
input [7:0] x2181 ,
input [7:0] x2182 ,
input [7:0] x2183 ,
input [7:0] x2184 ,
input [7:0] x2185 ,
input [7:0] x2186 ,
input [7:0] x2187 ,
input [7:0] x2188 ,
input [7:0] x2189 ,
input [7:0] x2190 ,
input [7:0] x2191 ,
input [7:0] x2192 ,
input [7:0] x2193 ,
input [7:0] x2194 ,
input [7:0] x2195 ,
input [7:0] x2196 ,
input [7:0] x2197 ,
input [7:0] x2198 ,
input [7:0] x2199 ,
input [7:0] x2200 ,
input [7:0] x2201 ,
input [7:0] x2202 ,
input [7:0] x2203 ,
input [7:0] x2204 ,
input [7:0] x2205 ,
input [7:0] x2206 ,
input [7:0] x2207 ,
input [7:0] x2208 ,
input [7:0] x2209 ,
input [7:0] x2210 ,
input [7:0] x2211 ,
input [7:0] x2212 ,
input [7:0] x2213 ,
input [7:0] x2214 ,
input [7:0] x2215 ,
input [7:0] x2216 ,
input [7:0] x2217 ,
input [7:0] x2218 ,
input [7:0] x2219 ,
input [7:0] x2220 ,
input [7:0] x2221 ,
input [7:0] x2222 ,
input [7:0] x2223 ,
input [7:0] x2224 ,
input [7:0] x2225 ,
input [7:0] x2226 ,
input [7:0] x2227 ,
input [7:0] x2228 ,
input [7:0] x2229 ,
input [7:0] x2230 ,
input [7:0] x2231 ,
input [7:0] x2232 ,
input [7:0] x2233 ,
input [7:0] x2234 ,
input [7:0] x2235 ,
input [7:0] x2236 ,
input [7:0] x2237 ,
input [7:0] x2238 ,
input [7:0] x2239 ,
input [7:0] x2240 ,
input [7:0] x2241 ,
input [7:0] x2242 ,
input [7:0] x2243 ,
input [7:0] x2244 ,
input [7:0] x2245 ,
input [7:0] x2246 ,
input [7:0] x2247 ,
input [7:0] x2248 ,
input [7:0] x2249 ,
input [7:0] x2250 ,
input [7:0] x2251 ,
input [7:0] x2252 ,
input [7:0] x2253 ,
input [7:0] x2254 ,
input [7:0] x2255 ,
input [7:0] x2256 ,
input [7:0] x2257 ,
input [7:0] x2258 ,
input [7:0] x2259 ,
input [7:0] x2260 ,
input [7:0] x2261 ,
input [7:0] x2262 ,
input [7:0] x2263 ,
input [7:0] x2264 ,
input [7:0] x2265 ,
input [7:0] x2266 ,
input [7:0] x2267 ,
input [7:0] x2268 ,
input [7:0] x2269 ,
input [7:0] x2270 ,
input [7:0] x2271 ,
input [7:0] x2272 ,
input [7:0] x2273 ,
input [7:0] x2274 ,
input [7:0] x2275 ,
input [7:0] x2276 ,
input [7:0] x2277 ,
input [7:0] x2278 ,
input [7:0] x2279 ,
input [7:0] x2280 ,
input [7:0] x2281 ,
input [7:0] x2282 ,
input [7:0] x2283 ,
input [7:0] x2284 ,
input [7:0] x2285 ,
input [7:0] x2286 ,
input [7:0] x2287 ,
input [7:0] x2288 ,
input [7:0] x2289 ,
input [7:0] x2290 ,
input [7:0] x2291 ,
input [7:0] x2292 ,
input [7:0] x2293 ,
input [7:0] x2294 ,
input [7:0] x2295 ,
input [7:0] x2296 ,
input [7:0] x2297 ,
input [7:0] x2298 ,
input [7:0] x2299 ,
input [7:0] x2300 ,
input [7:0] x2301 ,
input [7:0] x2302 ,
input [7:0] x2303 ,
input [7:0] x2304 ,
input [7:0] x2305 ,
input [7:0] x2306 ,
input [7:0] x2307 ,
input [7:0] x2308 ,
input [7:0] x2309 ,
input [7:0] x2310 ,
input [7:0] x2311 ,
input [7:0] x2312 ,
input [7:0] x2313 ,
input [7:0] x2314 ,
input [7:0] x2315 ,
input [7:0] x2316 ,
input [7:0] x2317 ,
input [7:0] x2318 ,
input [7:0] x2319 ,
input [7:0] x2320 ,
input [7:0] x2321 ,
input [7:0] x2322 ,
input [7:0] x2323 ,
input [7:0] x2324 ,
input [7:0] x2325 ,
input [7:0] x2326 ,
input [7:0] x2327 ,
input [7:0] x2328 ,
input [7:0] x2329 ,
input [7:0] x2330 ,
input [7:0] x2331 ,
input [7:0] x2332 ,
input [7:0] x2333 ,
input [7:0] x2334 ,
input [7:0] x2335 ,
input [7:0] x2336 ,
input [7:0] x2337 ,
input [7:0] x2338 ,
input [7:0] x2339 ,
input [7:0] x2340 ,
input [7:0] x2341 ,
input [7:0] x2342 ,
input [7:0] x2343 ,
input [7:0] x2344 ,
input [7:0] x2345 ,
input [7:0] x2346 ,
input [7:0] x2347 ,
input [7:0] x2348 ,
input [7:0] x2349 ,
input [7:0] x2350 ,
input [7:0] x2351 ,
input [7:0] x2352 ,
input [7:0] x2353 ,
input [7:0] x2354 ,
input [7:0] x2355 ,
input [7:0] x2356 ,
input [7:0] x2357 ,
input [7:0] x2358 ,
input [7:0] x2359 ,
input [7:0] x2360 ,
input [7:0] x2361 ,
input [7:0] x2362 ,
input [7:0] x2363 ,
input [7:0] x2364 ,
input [7:0] x2365 ,
input [7:0] x2366 ,
input [7:0] x2367 ,
input [7:0] x2368 ,
input [7:0] x2369 ,
input [7:0] x2370 ,
input [7:0] x2371 ,
input [7:0] x2372 ,
input [7:0] x2373 ,
input [7:0] x2374 ,
input [7:0] x2375 ,
input [7:0] x2376 ,
input [7:0] x2377 ,
input [7:0] x2378 ,
input [7:0] x2379 ,
input [7:0] x2380 ,
input [7:0] x2381 ,
input [7:0] x2382 ,
input [7:0] x2383 ,
input [7:0] x2384 ,
input [7:0] x2385 ,
input [7:0] x2386 ,
input [7:0] x2387 ,
input [7:0] x2388 ,
input [7:0] x2389 ,
input [7:0] x2390 ,
input [7:0] x2391 ,
input [7:0] x2392 ,
input [7:0] x2393 ,
input [7:0] x2394 ,
input [7:0] x2395 ,
input [7:0] x2396 ,
input [7:0] x2397 ,
input [7:0] x2398 ,
input [7:0] x2399 ,
input [7:0] x2400 ,
input [7:0] x2401 ,
input [7:0] x2402 ,
input [7:0] x2403 ,
input [7:0] x2404 ,
input [7:0] x2405 ,
input [7:0] x2406 ,
input [7:0] x2407 ,
input [7:0] x2408 ,
input [7:0] x2409 ,
input [7:0] x2410 ,
input [7:0] x2411 ,
input [7:0] x2412 ,
input [7:0] x2413 ,
input [7:0] x2414 ,
input [7:0] x2415 ,
input [7:0] x2416 ,
input [7:0] x2417 ,
input [7:0] x2418 ,
input [7:0] x2419 ,
input [7:0] x2420 ,
input [7:0] x2421 ,
input [7:0] x2422 ,
input [7:0] x2423 ,
input [7:0] x2424 ,
input [7:0] x2425 ,
input [7:0] x2426 ,
input [7:0] x2427 ,
input [7:0] x2428 ,
input [7:0] x2429 ,
input [7:0] x2430 ,
input [7:0] x2431 ,
input [7:0] x2432 ,
input [7:0] x2433 ,
input [7:0] x2434 ,
input [7:0] x2435 ,
input [7:0] x2436 ,
input [7:0] x2437 ,
input [7:0] x2438 ,
input [7:0] x2439 ,
input [7:0] x2440 ,
input [7:0] x2441 ,
input [7:0] x2442 ,
input [7:0] x2443 ,
input [7:0] x2444 ,
input [7:0] x2445 ,
input [7:0] x2446 ,
input [7:0] x2447 ,
input [7:0] x2448 ,
input [7:0] x2449 ,
input [7:0] x2450 ,
input [7:0] x2451 ,
input [7:0] x2452 ,
input [7:0] x2453 ,
input [7:0] x2454 ,
input [7:0] x2455 ,
input [7:0] x2456 ,
input [7:0] x2457 ,
input [7:0] x2458 ,
input [7:0] x2459 ,
input [7:0] x2460 ,
input [7:0] x2461 ,
input [7:0] x2462 ,
input [7:0] x2463 ,
input [7:0] x2464 ,
input [7:0] x2465 ,
input [7:0] x2466 ,
input [7:0] x2467 ,
input [7:0] x2468 ,
input [7:0] x2469 ,
input [7:0] x2470 ,
input [7:0] x2471 ,
input [7:0] x2472 ,
input [7:0] x2473 ,
input [7:0] x2474 ,
input [7:0] x2475 ,
input [7:0] x2476 ,
input [7:0] x2477 ,
input [7:0] x2478 ,
input [7:0] x2479 ,
input [7:0] x2480 ,
input [7:0] x2481 ,
input [7:0] x2482 ,
input [7:0] x2483 ,
input [7:0] x2484 ,
input [7:0] x2485 ,
input [7:0] x2486 ,
input [7:0] x2487 ,
input [7:0] x2488 ,
input [7:0] x2489 ,
input [7:0] x2490 ,
input [7:0] x2491 ,
input [7:0] x2492 ,
input [7:0] x2493 ,
input [7:0] x2494 ,
input [7:0] x2495 ,
input [7:0] x2496 ,
input [7:0] x2497 ,
input [7:0] x2498 ,
input [7:0] x2499 ,
input [7:0] x2500 ,
input [7:0] x2501 ,
input [7:0] x2502 ,
input [7:0] x2503 ,
input [7:0] x2504 ,
input [7:0] x2505 ,
input [7:0] x2506 ,
input [7:0] x2507 ,
input [7:0] x2508 ,
input [7:0] x2509 ,
input [7:0] x2510 ,
input [7:0] x2511 ,
input [7:0] x2512 ,
input [7:0] x2513 ,
input [7:0] x2514 ,
input [7:0] x2515 ,
input [7:0] x2516 ,
input [7:0] x2517 ,
input [7:0] x2518 ,
input [7:0] x2519 ,
input [7:0] x2520 ,
input [7:0] x2521 ,
input [7:0] x2522 ,
input [7:0] x2523 ,
input [7:0] x2524 ,
input [7:0] x2525 ,
input [7:0] x2526 ,
input [7:0] x2527 ,
input [7:0] x2528 ,
input [7:0] x2529 ,
input [7:0] x2530 ,
input [7:0] x2531 ,
input [7:0] x2532 ,
input [7:0] x2533 ,
input [7:0] x2534 ,
input [7:0] x2535 ,
input [7:0] x2536 ,
input [7:0] x2537 ,
input [7:0] x2538 ,
input [7:0] x2539 ,
input [7:0] x2540 ,
input [7:0] x2541 ,
input [7:0] x2542 ,
input [7:0] x2543 ,
input [7:0] x2544 ,
input [7:0] x2545 ,
input [7:0] x2546 ,
input [7:0] x2547 ,
input [7:0] x2548 ,
input [7:0] x2549 ,
input [7:0] x2550 ,
input [7:0] x2551 ,
input [7:0] x2552 ,
input [7:0] x2553 ,
input [7:0] x2554 ,
input [7:0] x2555 ,
input [7:0] x2556 ,
input [7:0] x2557 ,
input [7:0] x2558 ,
input [7:0] x2559 ,
input [7:0] x2560 ,
input [7:0] x2561 ,
input [7:0] x2562 ,
input [7:0] x2563 ,
input [7:0] x2564 ,
input [7:0] x2565 ,
input [7:0] x2566 ,
input [7:0] x2567 ,
input [7:0] x2568 ,
input [7:0] x2569 ,
input [7:0] x2570 ,
input [7:0] x2571 ,
input [7:0] x2572 ,
input [7:0] x2573 ,
input [7:0] x2574 ,
input [7:0] x2575 ,
input [7:0] x2576 ,
input [7:0] x2577 ,
input [7:0] x2578 ,
input [7:0] x2579 ,
input [7:0] x2580 ,
input [7:0] x2581 ,
input [7:0] x2582 ,
input [7:0] x2583 ,
input [7:0] x2584 ,
input [7:0] x2585 ,
input [7:0] x2586 ,
input [7:0] x2587 ,
input [7:0] x2588 ,
input [7:0] x2589 ,
input [7:0] x2590 ,
input [7:0] x2591 ,
input [7:0] x2592 ,
input [7:0] x2593 ,
input [7:0] x2594 ,
input [7:0] x2595 ,
input [7:0] x2596 ,
input [7:0] x2597 ,
input [7:0] x2598 ,
input [7:0] x2599 ,
input [7:0] x2600 ,
input [7:0] x2601 ,
input [7:0] x2602 ,
input [7:0] x2603 ,
input [7:0] x2604 ,
input [7:0] x2605 ,
input [7:0] x2606 ,
input [7:0] x2607 ,
input [7:0] x2608 ,
input [7:0] x2609 ,
input [7:0] x2610 ,
input [7:0] x2611 ,
input [7:0] x2612 ,
input [7:0] x2613 ,
input [7:0] x2614 ,
input [7:0] x2615 ,
input [7:0] x2616 ,
input [7:0] x2617 ,
input [7:0] x2618 ,
input [7:0] x2619 ,
input [7:0] x2620 ,
input [7:0] x2621 ,
input [7:0] x2622 ,
input [7:0] x2623 ,
input [7:0] x2624 ,
input [7:0] x2625 ,
input [7:0] x2626 ,
input [7:0] x2627 ,
input [7:0] x2628 ,
input [7:0] x2629 ,
input [7:0] x2630 ,
input [7:0] x2631 ,
input [7:0] x2632 ,
input [7:0] x2633 ,
input [7:0] x2634 ,
input [7:0] x2635 ,
input [7:0] x2636 ,
input [7:0] x2637 ,
input [7:0] x2638 ,
input [7:0] x2639 ,
input [7:0] x2640 ,
input [7:0] x2641 ,
input [7:0] x2642 ,
input [7:0] x2643 ,
input [7:0] x2644 ,
input [7:0] x2645 ,
input [7:0] x2646 ,
input [7:0] x2647 ,
input [7:0] x2648 ,
input [7:0] x2649 ,
input [7:0] x2650 ,
input [7:0] x2651 ,
input [7:0] x2652 ,
input [7:0] x2653 ,
input [7:0] x2654 ,
input [7:0] x2655 ,
input [7:0] x2656 ,
input [7:0] x2657 ,
input [7:0] x2658 ,
input [7:0] x2659 ,
input [7:0] x2660 ,
input [7:0] x2661 ,
input [7:0] x2662 ,
input [7:0] x2663 ,
input [7:0] x2664 ,
input [7:0] x2665 ,
input [7:0] x2666 ,
input [7:0] x2667 ,
input [7:0] x2668 ,
input [7:0] x2669 ,
input [7:0] x2670 ,
input [7:0] x2671 ,
input [7:0] x2672 ,
input [7:0] x2673 ,
input [7:0] x2674 ,
input [7:0] x2675 ,
input [7:0] x2676 ,
input [7:0] x2677 ,
input [7:0] x2678 ,
input [7:0] x2679 ,
input [7:0] x2680 ,
input [7:0] x2681 ,
input [7:0] x2682 ,
input [7:0] x2683 ,
input [7:0] x2684 ,
input [7:0] x2685 ,
input [7:0] x2686 ,
input [7:0] x2687 ,
input [7:0] x2688 ,
input [7:0] x2689 ,
input [7:0] x2690 ,
input [7:0] x2691 ,
input [7:0] x2692 ,
input [7:0] x2693 ,
input [7:0] x2694 ,
input [7:0] x2695 ,
input [7:0] x2696 ,
input [7:0] x2697 ,
input [7:0] x2698 ,
input [7:0] x2699 ,
input [7:0] x2700 ,
input [7:0] x2701 ,
input [7:0] x2702 ,
input [7:0] x2703 ,
input [7:0] x2704 ,
input [7:0] x2705 ,
input [7:0] x2706 ,
input [7:0] x2707 ,
input [7:0] x2708 ,
input [7:0] x2709 ,
input [7:0] x2710 ,
input [7:0] x2711 ,
input [7:0] x2712 ,
input [7:0] x2713 ,
input [7:0] x2714 ,
input [7:0] x2715 ,
input [7:0] x2716 ,
input [7:0] x2717 ,
input [7:0] x2718 ,
input [7:0] x2719 ,
input [7:0] x2720 ,
input [7:0] x2721 ,
input [7:0] x2722 ,
input [7:0] x2723 ,
input [7:0] x2724 ,
input [7:0] x2725 ,
input [7:0] x2726 ,
input [7:0] x2727 ,
input [7:0] x2728 ,
input [7:0] x2729 ,
input [7:0] x2730 ,
input [7:0] x2731 ,
input [7:0] x2732 ,
input [7:0] x2733 ,
input [7:0] x2734 ,
input [7:0] x2735 ,
input [7:0] x2736 ,
input [7:0] x2737 ,
input [7:0] x2738 ,
input [7:0] x2739 ,
input [7:0] x2740 ,
input [7:0] x2741 ,
input [7:0] x2742 ,
input [7:0] x2743 ,
input [7:0] x2744 ,
input [7:0] x2745 ,
input [7:0] x2746 ,
input [7:0] x2747 ,
input [7:0] x2748 ,
input [7:0] x2749 ,
input [7:0] x2750 ,
input [7:0] x2751 ,
input [7:0] x2752 ,
input [7:0] x2753 ,
input [7:0] x2754 ,
input [7:0] x2755 ,
input [7:0] x2756 ,
input [7:0] x2757 ,
input [7:0] x2758 ,
input [7:0] x2759 ,
input [7:0] x2760 ,
input [7:0] x2761 ,
input [7:0] x2762 ,
input [7:0] x2763 ,
input [7:0] x2764 ,
input [7:0] x2765 ,
input [7:0] x2766 ,
input [7:0] x2767 ,
input [7:0] x2768 ,
input [7:0] x2769 ,
input [7:0] x2770 ,
input [7:0] x2771 ,
input [7:0] x2772 ,
input [7:0] x2773 ,
input [7:0] x2774 ,
input [7:0] x2775 ,
input [7:0] x2776 ,
input [7:0] x2777 ,
input [7:0] x2778 ,
input [7:0] x2779 ,
input [7:0] x2780 ,
input [7:0] x2781 ,
input [7:0] x2782 ,
input [7:0] x2783 ,
input [7:0] x2784 ,
input [7:0] x2785 ,
input [7:0] x2786 ,
input [7:0] x2787 ,
input [7:0] x2788 ,
input [7:0] x2789 ,
input [7:0] x2790 ,
input [7:0] x2791 ,
input [7:0] x2792 ,
input [7:0] x2793 ,
input [7:0] x2794 ,
input [7:0] x2795 ,
input [7:0] x2796 ,
input [7:0] x2797 ,
input [7:0] x2798 ,
input [7:0] x2799 ,
input [7:0] x2800 ,
input [7:0] x2801 ,
input [7:0] x2802 ,
input [7:0] x2803 ,
input [7:0] x2804 ,
input [7:0] x2805 ,
input [7:0] x2806 ,
input [7:0] x2807 ,
input [7:0] x2808 ,
input [7:0] x2809 ,
input [7:0] x2810 ,
input [7:0] x2811 ,
input [7:0] x2812 ,
input [7:0] x2813 ,
input [7:0] x2814 ,
input [7:0] x2815 ,
input [7:0] x2816 ,
input [7:0] x2817 ,
input [7:0] x2818 ,
input [7:0] x2819 ,
input [7:0] x2820 ,
input [7:0] x2821 ,
input [7:0] x2822 ,
input [7:0] x2823 ,
input [7:0] x2824 ,
input [7:0] x2825 ,
input [7:0] x2826 ,
input [7:0] x2827 ,
input [7:0] x2828 ,
input [7:0] x2829 ,
input [7:0] x2830 ,
input [7:0] x2831 ,
input [7:0] x2832 ,
input [7:0] x2833 ,
input [7:0] x2834 ,
input [7:0] x2835 ,
input [7:0] x2836 ,
input [7:0] x2837 ,
input [7:0] x2838 ,
input [7:0] x2839 ,
input [7:0] x2840 ,
input [7:0] x2841 ,
input [7:0] x2842 ,
input [7:0] x2843 ,
input [7:0] x2844 ,
input [7:0] x2845 ,
input [7:0] x2846 ,
input [7:0] x2847 ,
input [7:0] x2848 ,
input [7:0] x2849 ,
input [7:0] x2850 ,
input [7:0] x2851 ,
input [7:0] x2852 ,
input [7:0] x2853 ,
input [7:0] x2854 ,
input [7:0] x2855 ,
input [7:0] x2856 ,
input [7:0] x2857 ,
input [7:0] x2858 ,
input [7:0] x2859 ,
input [7:0] x2860 ,
input [7:0] x2861 ,
input [7:0] x2862 ,
input [7:0] x2863 ,
input [7:0] x2864 ,
input [7:0] x2865 ,
input [7:0] x2866 ,
input [7:0] x2867 ,
input [7:0] x2868 ,
input [7:0] x2869 ,
input [7:0] x2870 ,
input [7:0] x2871 ,
input [7:0] x2872 ,
input [7:0] x2873 ,
input [7:0] x2874 ,
input [7:0] x2875 ,
input [7:0] x2876 ,
input [7:0] x2877 ,
input [7:0] x2878 ,
input [7:0] x2879 ,
input [7:0] x2880 ,
input [7:0] x2881 ,
input [7:0] x2882 ,
input [7:0] x2883 ,
input [7:0] x2884 ,
input [7:0] x2885 ,
input [7:0] x2886 ,
input [7:0] x2887 ,
input [7:0] x2888 ,
input [7:0] x2889 ,
input [7:0] x2890 ,
input [7:0] x2891 ,
input [7:0] x2892 ,
input [7:0] x2893 ,
input [7:0] x2894 ,
input [7:0] x2895 ,
input [7:0] x2896 ,
input [7:0] x2897 ,
input [7:0] x2898 ,
input [7:0] x2899 ,
input [7:0] x2900 ,
input [7:0] x2901 ,
input [7:0] x2902 ,
input [7:0] x2903 ,
input [7:0] x2904 ,
input [7:0] x2905 ,
input [7:0] x2906 ,
input [7:0] x2907 ,
input [7:0] x2908 ,
input [7:0] x2909 ,
input [7:0] x2910 ,
input [7:0] x2911 ,
input [7:0] x2912 ,
input [7:0] x2913 ,
input [7:0] x2914 ,
input [7:0] x2915 ,
input [7:0] x2916 ,
input [7:0] x2917 ,
input [7:0] x2918 ,
input [7:0] x2919 ,
input [7:0] x2920 ,
input [7:0] x2921 ,
input [7:0] x2922 ,
input [7:0] x2923 ,
input [7:0] x2924 ,
input [7:0] x2925 ,
input [7:0] x2926 ,
input [7:0] x2927 ,
input [7:0] x2928 ,
input [7:0] x2929 ,
input [7:0] x2930 ,
input [7:0] x2931 ,
input [7:0] x2932 ,
input [7:0] x2933 ,
input [7:0] x2934 ,
input [7:0] x2935 ,
input [7:0] x2936 ,
input [7:0] x2937 ,
input [7:0] x2938 ,
input [7:0] x2939 ,
input [7:0] x2940 ,
input [7:0] x2941 ,
input [7:0] x2942 ,
input [7:0] x2943 ,
input [7:0] x2944 ,
input [7:0] x2945 ,
input [7:0] x2946 ,
input [7:0] x2947 ,
input [7:0] x2948 ,
input [7:0] x2949 ,
input [7:0] x2950 ,
input [7:0] x2951 ,
input [7:0] x2952 ,
input [7:0] x2953 ,
input [7:0] x2954 ,
input [7:0] x2955 ,
input [7:0] x2956 ,
input [7:0] x2957 ,
input [7:0] x2958 ,
input [7:0] x2959 ,
input [7:0] x2960 ,
input [7:0] x2961 ,
input [7:0] x2962 ,
input [7:0] x2963 ,
input [7:0] x2964 ,
input [7:0] x2965 ,
input [7:0] x2966 ,
input [7:0] x2967 ,
input [7:0] x2968 ,
input [7:0] x2969 ,
input [7:0] x2970 ,
input [7:0] x2971 ,
input [7:0] x2972 ,
input [7:0] x2973 ,
input [7:0] x2974 ,
input [7:0] x2975 ,
input [7:0] x2976 ,
input [7:0] x2977 ,
input [7:0] x2978 ,
input [7:0] x2979 ,
input [7:0] x2980 ,
input [7:0] x2981 ,
input [7:0] x2982 ,
input [7:0] x2983 ,
input [7:0] x2984 ,
input [7:0] x2985 ,
input [7:0] x2986 ,
input [7:0] x2987 ,
input [7:0] x2988 ,
input [7:0] x2989 ,
input [7:0] x2990 ,
input [7:0] x2991 ,
input [7:0] x2992 ,
input [7:0] x2993 ,
input [7:0] x2994 ,
input [7:0] x2995 ,
input [7:0] x2996 ,
input [7:0] x2997 ,
input [7:0] x2998 ,
input [7:0] x2999 ,
input [7:0] x3000 ,
input [7:0] x3001 ,
input [7:0] x3002 ,
input [7:0] x3003 ,
input [7:0] x3004 ,
input [7:0] x3005 ,
input [7:0] x3006 ,
input [7:0] x3007 ,
input [7:0] x3008 ,
input [7:0] x3009 ,
input [7:0] x3010 ,
input [7:0] x3011 ,
input [7:0] x3012 ,
input [7:0] x3013 ,
input [7:0] x3014 ,
input [7:0] x3015 ,
input [7:0] x3016 ,
input [7:0] x3017 ,
input [7:0] x3018 ,
input [7:0] x3019 ,
input [7:0] x3020 ,
input [7:0] x3021 ,
input [7:0] x3022 ,
input [7:0] x3023 ,
input [7:0] x3024 ,
input [7:0] x3025 ,
input [7:0] x3026 ,
input [7:0] x3027 ,
input [7:0] x3028 ,
input [7:0] x3029 ,
input [7:0] x3030 ,
input [7:0] x3031 ,
input [7:0] x3032 ,
input [7:0] x3033 ,
input [7:0] x3034 ,
input [7:0] x3035 ,
input [7:0] x3036 ,
input [7:0] x3037 ,
input [7:0] x3038 ,
input [7:0] x3039 ,
input [7:0] x3040 ,
input [7:0] x3041 ,
input [7:0] x3042 ,
input [7:0] x3043 ,
input [7:0] x3044 ,
input [7:0] x3045 ,
input [7:0] x3046 ,
input [7:0] x3047 ,
input [7:0] x3048 ,
input [7:0] x3049 ,
input [7:0] x3050 ,
input [7:0] x3051 ,
input [7:0] x3052 ,
input [7:0] x3053 ,
input [7:0] x3054 ,
input [7:0] x3055 ,
input [7:0] x3056 ,
input [7:0] x3057 ,
input [7:0] x3058 ,
input [7:0] x3059 ,
input [7:0] x3060 ,
input [7:0] x3061 ,
input [7:0] x3062 ,
input [7:0] x3063 ,
input [7:0] x3064 ,
input [7:0] x3065 ,
input [7:0] x3066 ,
input [7:0] x3067 ,
input [7:0] x3068 ,
input [7:0] x3069 ,
input [7:0] x3070 ,
input [7:0] x3071 ,
output [6:0] y0 ,
output [6:0] y1 ,
output [6:0] y2 ,
output [6:0] y3 ,
output [6:0] y4 ,
output [6:0] y5 ,
output [6:0] y6 ,
output [6:0] y7 ,
output [6:0] y8 ,
output [6:0] y9 ,
output [6:0] y10 ,
output [6:0] y11 ,
output [6:0] y12 ,
output [6:0] y13 ,
output [6:0] y14 ,
output [6:0] y15 ,
output [6:0] y16 ,
output [6:0] y17 ,
output [6:0] y18 ,
output [6:0] y19 ,
output [6:0] y20 ,
output [6:0] y21 ,
output [6:0] y22 ,
output [6:0] y23 ,
output [6:0] y24 ,
output [6:0] y25 ,
output [6:0] y26 ,
output [6:0] y27 ,
output [6:0] y28 ,
output [6:0] y29 ,
output [6:0] y30 ,
output [6:0] y31 ,
output [6:0] y32 ,
output [6:0] y33 ,
output [6:0] y34 ,
output [6:0] y35 ,
output [6:0] y36 ,
output [6:0] y37 ,
output [6:0] y38 ,
output [6:0] y39 ,
output [6:0] y40 ,
output [6:0] y41 ,
output [6:0] y42 ,
output [6:0] y43 ,
output [6:0] y44 ,
output [6:0] y45 ,
output [6:0] y46 ,
output [6:0] y47 ,
output [6:0] y48 ,
output [6:0] y49 ,
output [6:0] y50 ,
output [6:0] y51 ,
output [6:0] y52 ,
output [6:0] y53 ,
output [6:0] y54 ,
output [6:0] y55 ,
output [6:0] y56 ,
output [6:0] y57 ,
output [6:0] y58 ,
output [6:0] y59 ,
output [6:0] y60 ,
output [6:0] y61 ,
output [6:0] y62 ,
output [6:0] y63 ,
output [6:0] y64 ,
output [6:0] y65 ,
output [6:0] y66 ,
output [6:0] y67 ,
output [6:0] y68 ,
output [6:0] y69 ,
output [6:0] y70 ,
output [6:0] y71 ,
output [6:0] y72 ,
output [6:0] y73 ,
output [6:0] y74 ,
output [6:0] y75 ,
output [6:0] y76 ,
output [6:0] y77 ,
output [6:0] y78 ,
output [6:0] y79 ,
output [6:0] y80 ,
output [6:0] y81 ,
output [6:0] y82 ,
output [6:0] y83 ,
output [6:0] y84 ,
output [6:0] y85 ,
output [6:0] y86 ,
output [6:0] y87 ,
output [6:0] y88 ,
output [6:0] y89 ,
output [6:0] y90 ,
output [6:0] y91 ,
output [6:0] y92 ,
output [6:0] y93 ,
output [6:0] y94 ,
output [6:0] y95 ,
output [6:0] y96 ,
output [6:0] y97 ,
output [6:0] y98 ,
output [6:0] y99 ,
output [6:0] y100 ,
output [6:0] y101 ,
output [6:0] y102 ,
output [6:0] y103 ,
output [6:0] y104 ,
output [6:0] y105 ,
output [6:0] y106 ,
output [6:0] y107 ,
output [6:0] y108 ,
output [6:0] y109 ,
output [6:0] y110 ,
output [6:0] y111 ,
output [6:0] y112 ,
output [6:0] y113 ,
output [6:0] y114 ,
output [6:0] y115 ,
output [6:0] y116 ,
output [6:0] y117 ,
output [6:0] y118 ,
output [6:0] y119 ,
output [6:0] y120 ,
output [6:0] y121 ,
output [6:0] y122 ,
output [6:0] y123 ,
output [6:0] y124 ,
output [6:0] y125 ,
output [6:0] y126 ,
output [6:0] y127 ,
output [6:0] y128 ,
output [6:0] y129 ,
output [6:0] y130 ,
output [6:0] y131 ,
output [6:0] y132 ,
output [6:0] y133 ,
output [6:0] y134 ,
output [6:0] y135 ,
output [6:0] y136 ,
output [6:0] y137 ,
output [6:0] y138 ,
output [6:0] y139 ,
output [6:0] y140 ,
output [6:0] y141 ,
output [6:0] y142 ,
output [6:0] y143 ,
output [6:0] y144 ,
output [6:0] y145 ,
output [6:0] y146 ,
output [6:0] y147 ,
output [6:0] y148 ,
output [6:0] y149 ,
output [6:0] y150 ,
output [6:0] y151 ,
output [6:0] y152 ,
output [6:0] y153 ,
output [6:0] y154 ,
output [6:0] y155 ,
output [6:0] y156 ,
output [6:0] y157 ,
output [6:0] y158 ,
output [6:0] y159 ,
output [6:0] y160 ,
output [6:0] y161 ,
output [6:0] y162 ,
output [6:0] y163 ,
output [6:0] y164 ,
output [6:0] y165 ,
output [6:0] y166 ,
output [6:0] y167 ,
output [6:0] y168 ,
output [6:0] y169 ,
output [6:0] y170 ,
output [6:0] y171 ,
output [6:0] y172 ,
output [6:0] y173 ,
output [6:0] y174 ,
output [6:0] y175 ,
output [6:0] y176 ,
output [6:0] y177 ,
output [6:0] y178 ,
output [6:0] y179 ,
output [6:0] y180 ,
output [6:0] y181 ,
output [6:0] y182 ,
output [6:0] y183 ,
output [6:0] y184 ,
output [6:0] y185 ,
output [6:0] y186 ,
output [6:0] y187 ,
output [6:0] y188 ,
output [6:0] y189 ,
output [6:0] y190 ,
output [6:0] y191 ,
output [6:0] y192 ,
output [6:0] y193 ,
output [6:0] y194 ,
output [6:0] y195 ,
output [6:0] y196 ,
output [6:0] y197 ,
output [6:0] y198 ,
output [6:0] y199 ,
output [6:0] y200 ,
output [6:0] y201 ,
output [6:0] y202 ,
output [6:0] y203 ,
output [6:0] y204 ,
output [6:0] y205 ,
output [6:0] y206 ,
output [6:0] y207 ,
output [6:0] y208 ,
output [6:0] y209 ,
output [6:0] y210 ,
output [6:0] y211 ,
output [6:0] y212 ,
output [6:0] y213 ,
output [6:0] y214 ,
output [6:0] y215 ,
output [6:0] y216 ,
output [6:0] y217 ,
output [6:0] y218 ,
output [6:0] y219 ,
output [6:0] y220 ,
output [6:0] y221 ,
output [6:0] y222 ,
output [6:0] y223 ,
output [6:0] y224 ,
output [6:0] y225 ,
output [6:0] y226 ,
output [6:0] y227 ,
output [6:0] y228 ,
output [6:0] y229 ,
output [6:0] y230 ,
output [6:0] y231 ,
output [6:0] y232 ,
output [6:0] y233 ,
output [6:0] y234 ,
output [6:0] y235 ,
output [6:0] y236 ,
output [6:0] y237 ,
output [6:0] y238 ,
output [6:0] y239 ,
output [6:0] y240 ,
output [6:0] y241 ,
output [6:0] y242 ,
output [6:0] y243 ,
output [6:0] y244 ,
output [6:0] y245 ,
output [6:0] y246 ,
output [6:0] y247 ,
output [6:0] y248 ,
output [6:0] y249 ,
output [6:0] y250 ,
output [6:0] y251 ,
output [6:0] y252 ,
output [6:0] y253 ,
output [6:0] y254 ,
output [6:0] y255 ,
output [6:0] y256 ,
output [6:0] y257 ,
output [6:0] y258 ,
output [6:0] y259 ,
output [6:0] y260 ,
output [6:0] y261 ,
output [6:0] y262 ,
output [6:0] y263 ,
output [6:0] y264 ,
output [6:0] y265 ,
output [6:0] y266 ,
output [6:0] y267 ,
output [6:0] y268 ,
output [6:0] y269 ,
output [6:0] y270 ,
output [6:0] y271 ,
output [6:0] y272 ,
output [6:0] y273 ,
output [6:0] y274 ,
output [6:0] y275 ,
output [6:0] y276 ,
output [6:0] y277 ,
output [6:0] y278 ,
output [6:0] y279 ,
output [6:0] y280 ,
output [6:0] y281 ,
output [6:0] y282 ,
output [6:0] y283 ,
output [6:0] y284 ,
output [6:0] y285 ,
output [6:0] y286 ,
output [6:0] y287 ,
output [6:0] y288 ,
output [6:0] y289 ,
output [6:0] y290 ,
output [6:0] y291 ,
output [6:0] y292 ,
output [6:0] y293 ,
output [6:0] y294 ,
output [6:0] y295 ,
output [6:0] y296 ,
output [6:0] y297 ,
output [6:0] y298 ,
output [6:0] y299 ,
output [6:0] y300 ,
output [6:0] y301 ,
output [6:0] y302 ,
output [6:0] y303 ,
output [6:0] y304 ,
output [6:0] y305 ,
output [6:0] y306 ,
output [6:0] y307 ,
output [6:0] y308 ,
output [6:0] y309 ,
output [6:0] y310 ,
output [6:0] y311 ,
output [6:0] y312 ,
output [6:0] y313 ,
output [6:0] y314 ,
output [6:0] y315 ,
output [6:0] y316 ,
output [6:0] y317 ,
output [6:0] y318 ,
output [6:0] y319 ,
output [6:0] y320 ,
output [6:0] y321 ,
output [6:0] y322 ,
output [6:0] y323 ,
output [6:0] y324 ,
output [6:0] y325 ,
output [6:0] y326 ,
output [6:0] y327 ,
output [6:0] y328 ,
output [6:0] y329 ,
output [6:0] y330 ,
output [6:0] y331 ,
output [6:0] y332 ,
output [6:0] y333 ,
output [6:0] y334 ,
output [6:0] y335 ,
output [6:0] y336 ,
output [6:0] y337 ,
output [6:0] y338 ,
output [6:0] y339 ,
output [6:0] y340 ,
output [6:0] y341 ,
output [6:0] y342 ,
output [6:0] y343 ,
output [6:0] y344 ,
output [6:0] y345 ,
output [6:0] y346 ,
output [6:0] y347 ,
output [6:0] y348 ,
output [6:0] y349 ,
output [6:0] y350 ,
output [6:0] y351 ,
output [6:0] y352 ,
output [6:0] y353 ,
output [6:0] y354 ,
output [6:0] y355 ,
output [6:0] y356 ,
output [6:0] y357 ,
output [6:0] y358 ,
output [6:0] y359 ,
output [6:0] y360 ,
output [6:0] y361 ,
output [6:0] y362 ,
output [6:0] y363 ,
output [6:0] y364 ,
output [6:0] y365 ,
output [6:0] y366 ,
output [6:0] y367 ,
output [6:0] y368 ,
output [6:0] y369 ,
output [6:0] y370 ,
output [6:0] y371 ,
output [6:0] y372 ,
output [6:0] y373 ,
output [6:0] y374 ,
output [6:0] y375 ,
output [6:0] y376 ,
output [6:0] y377 ,
output [6:0] y378 ,
output [6:0] y379 ,
output [6:0] y380 ,
output [6:0] y381 ,
output [6:0] y382 ,
output [6:0] y383 ,
output [6:0] y384 ,
output [6:0] y385 ,
output [6:0] y386 ,
output [6:0] y387 ,
output [6:0] y388 ,
output [6:0] y389 ,
output [6:0] y390 ,
output [6:0] y391 ,
output [6:0] y392 ,
output [6:0] y393 ,
output [6:0] y394 ,
output [6:0] y395 ,
output [6:0] y396 ,
output [6:0] y397 ,
output [6:0] y398 ,
output [6:0] y399 ,
output [6:0] y400 ,
output [6:0] y401 ,
output [6:0] y402 ,
output [6:0] y403 ,
output [6:0] y404 ,
output [6:0] y405 ,
output [6:0] y406 ,
output [6:0] y407 ,
output [6:0] y408 ,
output [6:0] y409 ,
output [6:0] y410 ,
output [6:0] y411 ,
output [6:0] y412 ,
output [6:0] y413 ,
output [6:0] y414 ,
output [6:0] y415 ,
output [6:0] y416 ,
output [6:0] y417 ,
output [6:0] y418 ,
output [6:0] y419 ,
output [6:0] y420 ,
output [6:0] y421 ,
output [6:0] y422 ,
output [6:0] y423 ,
output [6:0] y424 ,
output [6:0] y425 ,
output [6:0] y426 ,
output [6:0] y427 ,
output [6:0] y428 ,
output [6:0] y429 ,
output [6:0] y430 ,
output [6:0] y431 ,
output [6:0] y432 ,
output [6:0] y433 ,
output [6:0] y434 ,
output [6:0] y435 ,
output [6:0] y436 ,
output [6:0] y437 ,
output [6:0] y438 ,
output [6:0] y439 ,
output [6:0] y440 ,
output [6:0] y441 ,
output [6:0] y442 ,
output [6:0] y443 ,
output [6:0] y444 ,
output [6:0] y445 ,
output [6:0] y446 ,
output [6:0] y447 ,
output [6:0] y448 ,
output [6:0] y449 ,
output [6:0] y450 ,
output [6:0] y451 ,
output [6:0] y452 ,
output [6:0] y453 ,
output [6:0] y454 ,
output [6:0] y455 ,
output [6:0] y456 ,
output [6:0] y457 ,
output [6:0] y458 ,
output [6:0] y459 ,
output [6:0] y460 ,
output [6:0] y461 ,
output [6:0] y462 ,
output [6:0] y463 ,
output [6:0] y464 ,
output [6:0] y465 ,
output [6:0] y466 ,
output [6:0] y467 ,
output [6:0] y468 ,
output [6:0] y469 ,
output [6:0] y470 ,
output [6:0] y471 ,
output [6:0] y472 ,
output [6:0] y473 ,
output [6:0] y474 ,
output [6:0] y475 ,
output [6:0] y476 ,
output [6:0] y477 ,
output [6:0] y478 ,
output [6:0] y479 ,
output [6:0] y480 ,
output [6:0] y481 ,
output [6:0] y482 ,
output [6:0] y483 ,
output [6:0] y484 ,
output [6:0] y485 ,
output [6:0] y486 ,
output [6:0] y487 ,
output [6:0] y488 ,
output [6:0] y489 ,
output [6:0] y490 ,
output [6:0] y491 ,
output [6:0] y492 ,
output [6:0] y493 ,
output [6:0] y494 ,
output [6:0] y495 ,
output [6:0] y496 ,
output [6:0] y497 ,
output [6:0] y498 ,
output [6:0] y499 ,
output [6:0] y500 ,
output [6:0] y501 ,
output [6:0] y502 ,
output [6:0] y503 ,
output [6:0] y504 ,
output [6:0] y505 ,
output [6:0] y506 ,
output [6:0] y507 ,
output [6:0] y508 ,
output [6:0] y509 ,
output [6:0] y510 ,
output [6:0] y511 ,
output [6:0] y512 ,
output [6:0] y513 ,
output [6:0] y514 ,
output [6:0] y515 ,
output [6:0] y516 ,
output [6:0] y517 ,
output [6:0] y518 ,
output [6:0] y519 ,
output [6:0] y520 ,
output [6:0] y521 ,
output [6:0] y522 ,
output [6:0] y523 ,
output [6:0] y524 ,
output [6:0] y525 ,
output [6:0] y526 ,
output [6:0] y527 ,
output [6:0] y528 ,
output [6:0] y529 ,
output [6:0] y530 ,
output [6:0] y531 ,
output [6:0] y532 ,
output [6:0] y533 ,
output [6:0] y534 ,
output [6:0] y535 ,
output [6:0] y536 ,
output [6:0] y537 ,
output [6:0] y538 ,
output [6:0] y539 ,
output [6:0] y540 ,
output [6:0] y541 ,
output [6:0] y542 ,
output [6:0] y543 ,
output [6:0] y544 ,
output [6:0] y545 ,
output [6:0] y546 ,
output [6:0] y547 ,
output [6:0] y548 ,
output [6:0] y549 ,
output [6:0] y550 ,
output [6:0] y551 ,
output [6:0] y552 ,
output [6:0] y553 ,
output [6:0] y554 ,
output [6:0] y555 ,
output [6:0] y556 ,
output [6:0] y557 ,
output [6:0] y558 ,
output [6:0] y559 ,
output [6:0] y560 ,
output [6:0] y561 ,
output [6:0] y562 ,
output [6:0] y563 ,
output [6:0] y564 ,
output [6:0] y565 ,
output [6:0] y566 ,
output [6:0] y567 ,
output [6:0] y568 ,
output [6:0] y569 ,
output [6:0] y570 ,
output [6:0] y571 ,
output [6:0] y572 ,
output [6:0] y573 ,
output [6:0] y574 ,
output [6:0] y575 ,
output [6:0] y576 ,
output [6:0] y577 ,
output [6:0] y578 ,
output [6:0] y579 ,
output [6:0] y580 ,
output [6:0] y581 ,
output [6:0] y582 ,
output [6:0] y583 ,
output [6:0] y584 ,
output [6:0] y585 ,
output [6:0] y586 ,
output [6:0] y587 ,
output [6:0] y588 ,
output [6:0] y589 ,
output [6:0] y590 ,
output [6:0] y591 ,
output [6:0] y592 ,
output [6:0] y593 ,
output [6:0] y594 ,
output [6:0] y595 ,
output [6:0] y596 ,
output [6:0] y597 ,
output [6:0] y598 ,
output [6:0] y599 ,
output [6:0] y600 ,
output [6:0] y601 ,
output [6:0] y602 ,
output [6:0] y603 ,
output [6:0] y604 ,
output [6:0] y605 ,
output [6:0] y606 ,
output [6:0] y607 ,
output [6:0] y608 ,
output [6:0] y609 ,
output [6:0] y610 ,
output [6:0] y611 ,
output [6:0] y612 ,
output [6:0] y613 ,
output [6:0] y614 ,
output [6:0] y615 ,
output [6:0] y616 ,
output [6:0] y617 ,
output [6:0] y618 ,
output [6:0] y619 ,
output [6:0] y620 ,
output [6:0] y621 ,
output [6:0] y622 ,
output [6:0] y623 ,
output [6:0] y624 ,
output [6:0] y625 ,
output [6:0] y626 ,
output [6:0] y627 ,
output [6:0] y628 ,
output [6:0] y629 ,
output [6:0] y630 ,
output [6:0] y631 ,
output [6:0] y632 ,
output [6:0] y633 ,
output [6:0] y634 ,
output [6:0] y635 ,
output [6:0] y636 ,
output [6:0] y637 ,
output [6:0] y638 ,
output [6:0] y639 ,
output [6:0] y640 ,
output [6:0] y641 ,
output [6:0] y642 ,
output [6:0] y643 ,
output [6:0] y644 ,
output [6:0] y645 ,
output [6:0] y646 ,
output [6:0] y647 ,
output [6:0] y648 ,
output [6:0] y649 ,
output [6:0] y650 ,
output [6:0] y651 ,
output [6:0] y652 ,
output [6:0] y653 ,
output [6:0] y654 ,
output [6:0] y655 ,
output [6:0] y656 ,
output [6:0] y657 ,
output [6:0] y658 ,
output [6:0] y659 ,
output [6:0] y660 ,
output [6:0] y661 ,
output [6:0] y662 ,
output [6:0] y663 ,
output [6:0] y664 ,
output [6:0] y665 ,
output [6:0] y666 ,
output [6:0] y667 ,
output [6:0] y668 ,
output [6:0] y669 ,
output [6:0] y670 ,
output [6:0] y671 ,
output [6:0] y672 ,
output [6:0] y673 ,
output [6:0] y674 ,
output [6:0] y675 ,
output [6:0] y676 ,
output [6:0] y677 ,
output [6:0] y678 ,
output [6:0] y679 ,
output [6:0] y680 ,
output [6:0] y681 ,
output [6:0] y682 ,
output [6:0] y683 ,
output [6:0] y684 ,
output [6:0] y685 ,
output [6:0] y686 ,
output [6:0] y687 ,
output [6:0] y688 ,
output [6:0] y689 ,
output [6:0] y690 ,
output [6:0] y691 ,
output [6:0] y692 ,
output [6:0] y693 ,
output [6:0] y694 ,
output [6:0] y695 ,
output [6:0] y696 ,
output [6:0] y697 ,
output [6:0] y698 ,
output [6:0] y699 ,
output [6:0] y700 ,
output [6:0] y701 ,
output [6:0] y702 ,
output [6:0] y703 ,
output [6:0] y704 ,
output [6:0] y705 ,
output [6:0] y706 ,
output [6:0] y707 ,
output [6:0] y708 ,
output [6:0] y709 ,
output [6:0] y710 ,
output [6:0] y711 ,
output [6:0] y712 ,
output [6:0] y713 ,
output [6:0] y714 ,
output [6:0] y715 ,
output [6:0] y716 ,
output [6:0] y717 ,
output [6:0] y718 ,
output [6:0] y719 ,
output [6:0] y720 ,
output [6:0] y721 ,
output [6:0] y722 ,
output [6:0] y723 ,
output [6:0] y724 ,
output [6:0] y725 ,
output [6:0] y726 ,
output [6:0] y727 ,
output [6:0] y728 ,
output [6:0] y729 ,
output [6:0] y730 ,
output [6:0] y731 ,
output [6:0] y732 ,
output [6:0] y733 ,
output [6:0] y734 ,
output [6:0] y735 ,
output [6:0] y736 ,
output [6:0] y737 ,
output [6:0] y738 ,
output [6:0] y739 ,
output [6:0] y740 ,
output [6:0] y741 ,
output [6:0] y742 ,
output [6:0] y743 ,
output [6:0] y744 ,
output [6:0] y745 ,
output [6:0] y746 ,
output [6:0] y747 ,
output [6:0] y748 ,
output [6:0] y749 ,
output [6:0] y750 ,
output [6:0] y751 ,
output [6:0] y752 ,
output [6:0] y753 ,
output [6:0] y754 ,
output [6:0] y755 ,
output [6:0] y756 ,
output [6:0] y757 ,
output [6:0] y758 ,
output [6:0] y759 ,
output [6:0] y760 ,
output [6:0] y761 ,
output [6:0] y762 ,
output [6:0] y763 ,
output [6:0] y764 ,
output [6:0] y765 ,
output [6:0] y766 ,
output [6:0] y767 
);
assign y0=x0[7:1];
assign y256=x1024[7:1];
assign y512=x2048[7:1];
assign y1=x2[7:1];
assign y257=x1026[7:1];
assign y513=x2050[7:1];
assign y2=x4[7:1];
assign y258=x1028[7:1];
assign y514=x2052[7:1];
assign y3=x6[7:1];
assign y259=x1030[7:1];
assign y515=x2054[7:1];
assign y4=x8[7:1];
assign y260=x1032[7:1];
assign y516=x2056[7:1];
assign y5=x10[7:1];
assign y261=x1034[7:1];
assign y517=x2058[7:1];
assign y6=x12[7:1];
assign y262=x1036[7:1];
assign y518=x2060[7:1];
assign y7=x14[7:1];
assign y263=x1038[7:1];
assign y519=x2062[7:1];
assign y8=x16[7:1];
assign y264=x1040[7:1];
assign y520=x2064[7:1];
assign y9=x18[7:1];
assign y265=x1042[7:1];
assign y521=x2066[7:1];
assign y10=x20[7:1];
assign y266=x1044[7:1];
assign y522=x2068[7:1];
assign y11=x22[7:1];
assign y267=x1046[7:1];
assign y523=x2070[7:1];
assign y12=x24[7:1];
assign y268=x1048[7:1];
assign y524=x2072[7:1];
assign y13=x26[7:1];
assign y269=x1050[7:1];
assign y525=x2074[7:1];
assign y14=x28[7:1];
assign y270=x1052[7:1];
assign y526=x2076[7:1];
assign y15=x30[7:1];
assign y271=x1054[7:1];
assign y527=x2078[7:1];
assign y16=x64[7:1];
assign y272=x1088[7:1];
assign y528=x2112[7:1];
assign y17=x66[7:1];
assign y273=x1090[7:1];
assign y529=x2114[7:1];
assign y18=x68[7:1];
assign y274=x1092[7:1];
assign y530=x2116[7:1];
assign y19=x70[7:1];
assign y275=x1094[7:1];
assign y531=x2118[7:1];
assign y20=x72[7:1];
assign y276=x1096[7:1];
assign y532=x2120[7:1];
assign y21=x74[7:1];
assign y277=x1098[7:1];
assign y533=x2122[7:1];
assign y22=x76[7:1];
assign y278=x1100[7:1];
assign y534=x2124[7:1];
assign y23=x78[7:1];
assign y279=x1102[7:1];
assign y535=x2126[7:1];
assign y24=x80[7:1];
assign y280=x1104[7:1];
assign y536=x2128[7:1];
assign y25=x82[7:1];
assign y281=x1106[7:1];
assign y537=x2130[7:1];
assign y26=x84[7:1];
assign y282=x1108[7:1];
assign y538=x2132[7:1];
assign y27=x86[7:1];
assign y283=x1110[7:1];
assign y539=x2134[7:1];
assign y28=x88[7:1];
assign y284=x1112[7:1];
assign y540=x2136[7:1];
assign y29=x90[7:1];
assign y285=x1114[7:1];
assign y541=x2138[7:1];
assign y30=x92[7:1];
assign y286=x1116[7:1];
assign y542=x2140[7:1];
assign y31=x94[7:1];
assign y287=x1118[7:1];
assign y543=x2142[7:1];
assign y32=x128[7:1];
assign y288=x1152[7:1];
assign y544=x2176[7:1];
assign y33=x130[7:1];
assign y289=x1154[7:1];
assign y545=x2178[7:1];
assign y34=x132[7:1];
assign y290=x1156[7:1];
assign y546=x2180[7:1];
assign y35=x134[7:1];
assign y291=x1158[7:1];
assign y547=x2182[7:1];
assign y36=x136[7:1];
assign y292=x1160[7:1];
assign y548=x2184[7:1];
assign y37=x138[7:1];
assign y293=x1162[7:1];
assign y549=x2186[7:1];
assign y38=x140[7:1];
assign y294=x1164[7:1];
assign y550=x2188[7:1];
assign y39=x142[7:1];
assign y295=x1166[7:1];
assign y551=x2190[7:1];
assign y40=x144[7:1];
assign y296=x1168[7:1];
assign y552=x2192[7:1];
assign y41=x146[7:1];
assign y297=x1170[7:1];
assign y553=x2194[7:1];
assign y42=x148[7:1];
assign y298=x1172[7:1];
assign y554=x2196[7:1];
assign y43=x150[7:1];
assign y299=x1174[7:1];
assign y555=x2198[7:1];
assign y44=x152[7:1];
assign y300=x1176[7:1];
assign y556=x2200[7:1];
assign y45=x154[7:1];
assign y301=x1178[7:1];
assign y557=x2202[7:1];
assign y46=x156[7:1];
assign y302=x1180[7:1];
assign y558=x2204[7:1];
assign y47=x158[7:1];
assign y303=x1182[7:1];
assign y559=x2206[7:1];
assign y48=x192[7:1];
assign y304=x1216[7:1];
assign y560=x2240[7:1];
assign y49=x194[7:1];
assign y305=x1218[7:1];
assign y561=x2242[7:1];
assign y50=x196[7:1];
assign y306=x1220[7:1];
assign y562=x2244[7:1];
assign y51=x198[7:1];
assign y307=x1222[7:1];
assign y563=x2246[7:1];
assign y52=x200[7:1];
assign y308=x1224[7:1];
assign y564=x2248[7:1];
assign y53=x202[7:1];
assign y309=x1226[7:1];
assign y565=x2250[7:1];
assign y54=x204[7:1];
assign y310=x1228[7:1];
assign y566=x2252[7:1];
assign y55=x206[7:1];
assign y311=x1230[7:1];
assign y567=x2254[7:1];
assign y56=x208[7:1];
assign y312=x1232[7:1];
assign y568=x2256[7:1];
assign y57=x210[7:1];
assign y313=x1234[7:1];
assign y569=x2258[7:1];
assign y58=x212[7:1];
assign y314=x1236[7:1];
assign y570=x2260[7:1];
assign y59=x214[7:1];
assign y315=x1238[7:1];
assign y571=x2262[7:1];
assign y60=x216[7:1];
assign y316=x1240[7:1];
assign y572=x2264[7:1];
assign y61=x218[7:1];
assign y317=x1242[7:1];
assign y573=x2266[7:1];
assign y62=x220[7:1];
assign y318=x1244[7:1];
assign y574=x2268[7:1];
assign y63=x222[7:1];
assign y319=x1246[7:1];
assign y575=x2270[7:1];
assign y64=x256[7:1];
assign y320=x1280[7:1];
assign y576=x2304[7:1];
assign y65=x258[7:1];
assign y321=x1282[7:1];
assign y577=x2306[7:1];
assign y66=x260[7:1];
assign y322=x1284[7:1];
assign y578=x2308[7:1];
assign y67=x262[7:1];
assign y323=x1286[7:1];
assign y579=x2310[7:1];
assign y68=x264[7:1];
assign y324=x1288[7:1];
assign y580=x2312[7:1];
assign y69=x266[7:1];
assign y325=x1290[7:1];
assign y581=x2314[7:1];
assign y70=x268[7:1];
assign y326=x1292[7:1];
assign y582=x2316[7:1];
assign y71=x270[7:1];
assign y327=x1294[7:1];
assign y583=x2318[7:1];
assign y72=x272[7:1];
assign y328=x1296[7:1];
assign y584=x2320[7:1];
assign y73=x274[7:1];
assign y329=x1298[7:1];
assign y585=x2322[7:1];
assign y74=x276[7:1];
assign y330=x1300[7:1];
assign y586=x2324[7:1];
assign y75=x278[7:1];
assign y331=x1302[7:1];
assign y587=x2326[7:1];
assign y76=x280[7:1];
assign y332=x1304[7:1];
assign y588=x2328[7:1];
assign y77=x282[7:1];
assign y333=x1306[7:1];
assign y589=x2330[7:1];
assign y78=x284[7:1];
assign y334=x1308[7:1];
assign y590=x2332[7:1];
assign y79=x286[7:1];
assign y335=x1310[7:1];
assign y591=x2334[7:1];
assign y80=x320[7:1];
assign y336=x1344[7:1];
assign y592=x2368[7:1];
assign y81=x322[7:1];
assign y337=x1346[7:1];
assign y593=x2370[7:1];
assign y82=x324[7:1];
assign y338=x1348[7:1];
assign y594=x2372[7:1];
assign y83=x326[7:1];
assign y339=x1350[7:1];
assign y595=x2374[7:1];
assign y84=x328[7:1];
assign y340=x1352[7:1];
assign y596=x2376[7:1];
assign y85=x330[7:1];
assign y341=x1354[7:1];
assign y597=x2378[7:1];
assign y86=x332[7:1];
assign y342=x1356[7:1];
assign y598=x2380[7:1];
assign y87=x334[7:1];
assign y343=x1358[7:1];
assign y599=x2382[7:1];
assign y88=x336[7:1];
assign y344=x1360[7:1];
assign y600=x2384[7:1];
assign y89=x338[7:1];
assign y345=x1362[7:1];
assign y601=x2386[7:1];
assign y90=x340[7:1];
assign y346=x1364[7:1];
assign y602=x2388[7:1];
assign y91=x342[7:1];
assign y347=x1366[7:1];
assign y603=x2390[7:1];
assign y92=x344[7:1];
assign y348=x1368[7:1];
assign y604=x2392[7:1];
assign y93=x346[7:1];
assign y349=x1370[7:1];
assign y605=x2394[7:1];
assign y94=x348[7:1];
assign y350=x1372[7:1];
assign y606=x2396[7:1];
assign y95=x350[7:1];
assign y351=x1374[7:1];
assign y607=x2398[7:1];
assign y96=x384[7:1];
assign y352=x1408[7:1];
assign y608=x2432[7:1];
assign y97=x386[7:1];
assign y353=x1410[7:1];
assign y609=x2434[7:1];
assign y98=x388[7:1];
assign y354=x1412[7:1];
assign y610=x2436[7:1];
assign y99=x390[7:1];
assign y355=x1414[7:1];
assign y611=x2438[7:1];
assign y100=x392[7:1];
assign y356=x1416[7:1];
assign y612=x2440[7:1];
assign y101=x394[7:1];
assign y357=x1418[7:1];
assign y613=x2442[7:1];
assign y102=x396[7:1];
assign y358=x1420[7:1];
assign y614=x2444[7:1];
assign y103=x398[7:1];
assign y359=x1422[7:1];
assign y615=x2446[7:1];
assign y104=x400[7:1];
assign y360=x1424[7:1];
assign y616=x2448[7:1];
assign y105=x402[7:1];
assign y361=x1426[7:1];
assign y617=x2450[7:1];
assign y106=x404[7:1];
assign y362=x1428[7:1];
assign y618=x2452[7:1];
assign y107=x406[7:1];
assign y363=x1430[7:1];
assign y619=x2454[7:1];
assign y108=x408[7:1];
assign y364=x1432[7:1];
assign y620=x2456[7:1];
assign y109=x410[7:1];
assign y365=x1434[7:1];
assign y621=x2458[7:1];
assign y110=x412[7:1];
assign y366=x1436[7:1];
assign y622=x2460[7:1];
assign y111=x414[7:1];
assign y367=x1438[7:1];
assign y623=x2462[7:1];
assign y112=x448[7:1];
assign y368=x1472[7:1];
assign y624=x2496[7:1];
assign y113=x450[7:1];
assign y369=x1474[7:1];
assign y625=x2498[7:1];
assign y114=x452[7:1];
assign y370=x1476[7:1];
assign y626=x2500[7:1];
assign y115=x454[7:1];
assign y371=x1478[7:1];
assign y627=x2502[7:1];
assign y116=x456[7:1];
assign y372=x1480[7:1];
assign y628=x2504[7:1];
assign y117=x458[7:1];
assign y373=x1482[7:1];
assign y629=x2506[7:1];
assign y118=x460[7:1];
assign y374=x1484[7:1];
assign y630=x2508[7:1];
assign y119=x462[7:1];
assign y375=x1486[7:1];
assign y631=x2510[7:1];
assign y120=x464[7:1];
assign y376=x1488[7:1];
assign y632=x2512[7:1];
assign y121=x466[7:1];
assign y377=x1490[7:1];
assign y633=x2514[7:1];
assign y122=x468[7:1];
assign y378=x1492[7:1];
assign y634=x2516[7:1];
assign y123=x470[7:1];
assign y379=x1494[7:1];
assign y635=x2518[7:1];
assign y124=x472[7:1];
assign y380=x1496[7:1];
assign y636=x2520[7:1];
assign y125=x474[7:1];
assign y381=x1498[7:1];
assign y637=x2522[7:1];
assign y126=x476[7:1];
assign y382=x1500[7:1];
assign y638=x2524[7:1];
assign y127=x478[7:1];
assign y383=x1502[7:1];
assign y639=x2526[7:1];
assign y128=x512[7:1];
assign y384=x1536[7:1];
assign y640=x2560[7:1];
assign y129=x514[7:1];
assign y385=x1538[7:1];
assign y641=x2562[7:1];
assign y130=x516[7:1];
assign y386=x1540[7:1];
assign y642=x2564[7:1];
assign y131=x518[7:1];
assign y387=x1542[7:1];
assign y643=x2566[7:1];
assign y132=x520[7:1];
assign y388=x1544[7:1];
assign y644=x2568[7:1];
assign y133=x522[7:1];
assign y389=x1546[7:1];
assign y645=x2570[7:1];
assign y134=x524[7:1];
assign y390=x1548[7:1];
assign y646=x2572[7:1];
assign y135=x526[7:1];
assign y391=x1550[7:1];
assign y647=x2574[7:1];
assign y136=x528[7:1];
assign y392=x1552[7:1];
assign y648=x2576[7:1];
assign y137=x530[7:1];
assign y393=x1554[7:1];
assign y649=x2578[7:1];
assign y138=x532[7:1];
assign y394=x1556[7:1];
assign y650=x2580[7:1];
assign y139=x534[7:1];
assign y395=x1558[7:1];
assign y651=x2582[7:1];
assign y140=x536[7:1];
assign y396=x1560[7:1];
assign y652=x2584[7:1];
assign y141=x538[7:1];
assign y397=x1562[7:1];
assign y653=x2586[7:1];
assign y142=x540[7:1];
assign y398=x1564[7:1];
assign y654=x2588[7:1];
assign y143=x542[7:1];
assign y399=x1566[7:1];
assign y655=x2590[7:1];
assign y144=x576[7:1];
assign y400=x1600[7:1];
assign y656=x2624[7:1];
assign y145=x578[7:1];
assign y401=x1602[7:1];
assign y657=x2626[7:1];
assign y146=x580[7:1];
assign y402=x1604[7:1];
assign y658=x2628[7:1];
assign y147=x582[7:1];
assign y403=x1606[7:1];
assign y659=x2630[7:1];
assign y148=x584[7:1];
assign y404=x1608[7:1];
assign y660=x2632[7:1];
assign y149=x586[7:1];
assign y405=x1610[7:1];
assign y661=x2634[7:1];
assign y150=x588[7:1];
assign y406=x1612[7:1];
assign y662=x2636[7:1];
assign y151=x590[7:1];
assign y407=x1614[7:1];
assign y663=x2638[7:1];
assign y152=x592[7:1];
assign y408=x1616[7:1];
assign y664=x2640[7:1];
assign y153=x594[7:1];
assign y409=x1618[7:1];
assign y665=x2642[7:1];
assign y154=x596[7:1];
assign y410=x1620[7:1];
assign y666=x2644[7:1];
assign y155=x598[7:1];
assign y411=x1622[7:1];
assign y667=x2646[7:1];
assign y156=x600[7:1];
assign y412=x1624[7:1];
assign y668=x2648[7:1];
assign y157=x602[7:1];
assign y413=x1626[7:1];
assign y669=x2650[7:1];
assign y158=x604[7:1];
assign y414=x1628[7:1];
assign y670=x2652[7:1];
assign y159=x606[7:1];
assign y415=x1630[7:1];
assign y671=x2654[7:1];
assign y160=x640[7:1];
assign y416=x1664[7:1];
assign y672=x2688[7:1];
assign y161=x642[7:1];
assign y417=x1666[7:1];
assign y673=x2690[7:1];
assign y162=x644[7:1];
assign y418=x1668[7:1];
assign y674=x2692[7:1];
assign y163=x646[7:1];
assign y419=x1670[7:1];
assign y675=x2694[7:1];
assign y164=x648[7:1];
assign y420=x1672[7:1];
assign y676=x2696[7:1];
assign y165=x650[7:1];
assign y421=x1674[7:1];
assign y677=x2698[7:1];
assign y166=x652[7:1];
assign y422=x1676[7:1];
assign y678=x2700[7:1];
assign y167=x654[7:1];
assign y423=x1678[7:1];
assign y679=x2702[7:1];
assign y168=x656[7:1];
assign y424=x1680[7:1];
assign y680=x2704[7:1];
assign y169=x658[7:1];
assign y425=x1682[7:1];
assign y681=x2706[7:1];
assign y170=x660[7:1];
assign y426=x1684[7:1];
assign y682=x2708[7:1];
assign y171=x662[7:1];
assign y427=x1686[7:1];
assign y683=x2710[7:1];
assign y172=x664[7:1];
assign y428=x1688[7:1];
assign y684=x2712[7:1];
assign y173=x666[7:1];
assign y429=x1690[7:1];
assign y685=x2714[7:1];
assign y174=x668[7:1];
assign y430=x1692[7:1];
assign y686=x2716[7:1];
assign y175=x670[7:1];
assign y431=x1694[7:1];
assign y687=x2718[7:1];
assign y176=x704[7:1];
assign y432=x1728[7:1];
assign y688=x2752[7:1];
assign y177=x706[7:1];
assign y433=x1730[7:1];
assign y689=x2754[7:1];
assign y178=x708[7:1];
assign y434=x1732[7:1];
assign y690=x2756[7:1];
assign y179=x710[7:1];
assign y435=x1734[7:1];
assign y691=x2758[7:1];
assign y180=x712[7:1];
assign y436=x1736[7:1];
assign y692=x2760[7:1];
assign y181=x714[7:1];
assign y437=x1738[7:1];
assign y693=x2762[7:1];
assign y182=x716[7:1];
assign y438=x1740[7:1];
assign y694=x2764[7:1];
assign y183=x718[7:1];
assign y439=x1742[7:1];
assign y695=x2766[7:1];
assign y184=x720[7:1];
assign y440=x1744[7:1];
assign y696=x2768[7:1];
assign y185=x722[7:1];
assign y441=x1746[7:1];
assign y697=x2770[7:1];
assign y186=x724[7:1];
assign y442=x1748[7:1];
assign y698=x2772[7:1];
assign y187=x726[7:1];
assign y443=x1750[7:1];
assign y699=x2774[7:1];
assign y188=x728[7:1];
assign y444=x1752[7:1];
assign y700=x2776[7:1];
assign y189=x730[7:1];
assign y445=x1754[7:1];
assign y701=x2778[7:1];
assign y190=x732[7:1];
assign y446=x1756[7:1];
assign y702=x2780[7:1];
assign y191=x734[7:1];
assign y447=x1758[7:1];
assign y703=x2782[7:1];
assign y192=x768[7:1];
assign y448=x1792[7:1];
assign y704=x2816[7:1];
assign y193=x770[7:1];
assign y449=x1794[7:1];
assign y705=x2818[7:1];
assign y194=x772[7:1];
assign y450=x1796[7:1];
assign y706=x2820[7:1];
assign y195=x774[7:1];
assign y451=x1798[7:1];
assign y707=x2822[7:1];
assign y196=x776[7:1];
assign y452=x1800[7:1];
assign y708=x2824[7:1];
assign y197=x778[7:1];
assign y453=x1802[7:1];
assign y709=x2826[7:1];
assign y198=x780[7:1];
assign y454=x1804[7:1];
assign y710=x2828[7:1];
assign y199=x782[7:1];
assign y455=x1806[7:1];
assign y711=x2830[7:1];
assign y200=x784[7:1];
assign y456=x1808[7:1];
assign y712=x2832[7:1];
assign y201=x786[7:1];
assign y457=x1810[7:1];
assign y713=x2834[7:1];
assign y202=x788[7:1];
assign y458=x1812[7:1];
assign y714=x2836[7:1];
assign y203=x790[7:1];
assign y459=x1814[7:1];
assign y715=x2838[7:1];
assign y204=x792[7:1];
assign y460=x1816[7:1];
assign y716=x2840[7:1];
assign y205=x794[7:1];
assign y461=x1818[7:1];
assign y717=x2842[7:1];
assign y206=x796[7:1];
assign y462=x1820[7:1];
assign y718=x2844[7:1];
assign y207=x798[7:1];
assign y463=x1822[7:1];
assign y719=x2846[7:1];
assign y208=x832[7:1];
assign y464=x1856[7:1];
assign y720=x2880[7:1];
assign y209=x834[7:1];
assign y465=x1858[7:1];
assign y721=x2882[7:1];
assign y210=x836[7:1];
assign y466=x1860[7:1];
assign y722=x2884[7:1];
assign y211=x838[7:1];
assign y467=x1862[7:1];
assign y723=x2886[7:1];
assign y212=x840[7:1];
assign y468=x1864[7:1];
assign y724=x2888[7:1];
assign y213=x842[7:1];
assign y469=x1866[7:1];
assign y725=x2890[7:1];
assign y214=x844[7:1];
assign y470=x1868[7:1];
assign y726=x2892[7:1];
assign y215=x846[7:1];
assign y471=x1870[7:1];
assign y727=x2894[7:1];
assign y216=x848[7:1];
assign y472=x1872[7:1];
assign y728=x2896[7:1];
assign y217=x850[7:1];
assign y473=x1874[7:1];
assign y729=x2898[7:1];
assign y218=x852[7:1];
assign y474=x1876[7:1];
assign y730=x2900[7:1];
assign y219=x854[7:1];
assign y475=x1878[7:1];
assign y731=x2902[7:1];
assign y220=x856[7:1];
assign y476=x1880[7:1];
assign y732=x2904[7:1];
assign y221=x858[7:1];
assign y477=x1882[7:1];
assign y733=x2906[7:1];
assign y222=x860[7:1];
assign y478=x1884[7:1];
assign y734=x2908[7:1];
assign y223=x862[7:1];
assign y479=x1886[7:1];
assign y735=x2910[7:1];
assign y224=x896[7:1];
assign y480=x1920[7:1];
assign y736=x2944[7:1];
assign y225=x898[7:1];
assign y481=x1922[7:1];
assign y737=x2946[7:1];
assign y226=x900[7:1];
assign y482=x1924[7:1];
assign y738=x2948[7:1];
assign y227=x902[7:1];
assign y483=x1926[7:1];
assign y739=x2950[7:1];
assign y228=x904[7:1];
assign y484=x1928[7:1];
assign y740=x2952[7:1];
assign y229=x906[7:1];
assign y485=x1930[7:1];
assign y741=x2954[7:1];
assign y230=x908[7:1];
assign y486=x1932[7:1];
assign y742=x2956[7:1];
assign y231=x910[7:1];
assign y487=x1934[7:1];
assign y743=x2958[7:1];
assign y232=x912[7:1];
assign y488=x1936[7:1];
assign y744=x2960[7:1];
assign y233=x914[7:1];
assign y489=x1938[7:1];
assign y745=x2962[7:1];
assign y234=x916[7:1];
assign y490=x1940[7:1];
assign y746=x2964[7:1];
assign y235=x918[7:1];
assign y491=x1942[7:1];
assign y747=x2966[7:1];
assign y236=x920[7:1];
assign y492=x1944[7:1];
assign y748=x2968[7:1];
assign y237=x922[7:1];
assign y493=x1946[7:1];
assign y749=x2970[7:1];
assign y238=x924[7:1];
assign y494=x1948[7:1];
assign y750=x2972[7:1];
assign y239=x926[7:1];
assign y495=x1950[7:1];
assign y751=x2974[7:1];
assign y240=x960[7:1];
assign y496=x1984[7:1];
assign y752=x3008[7:1];
assign y241=x962[7:1];
assign y497=x1986[7:1];
assign y753=x3010[7:1];
assign y242=x964[7:1];
assign y498=x1988[7:1];
assign y754=x3012[7:1];
assign y243=x966[7:1];
assign y499=x1990[7:1];
assign y755=x3014[7:1];
assign y244=x968[7:1];
assign y500=x1992[7:1];
assign y756=x3016[7:1];
assign y245=x970[7:1];
assign y501=x1994[7:1];
assign y757=x3018[7:1];
assign y246=x972[7:1];
assign y502=x1996[7:1];
assign y758=x3020[7:1];
assign y247=x974[7:1];
assign y503=x1998[7:1];
assign y759=x3022[7:1];
assign y248=x976[7:1];
assign y504=x2000[7:1];
assign y760=x3024[7:1];
assign y249=x978[7:1];
assign y505=x2002[7:1];
assign y761=x3026[7:1];
assign y250=x980[7:1];
assign y506=x2004[7:1];
assign y762=x3028[7:1];
assign y251=x982[7:1];
assign y507=x2006[7:1];
assign y763=x3030[7:1];
assign y252=x984[7:1];
assign y508=x2008[7:1];
assign y764=x3032[7:1];
assign y253=x986[7:1];
assign y509=x2010[7:1];
assign y765=x3034[7:1];
assign y254=x988[7:1];
assign y510=x2012[7:1];
assign y766=x3036[7:1];
assign y255=x990[7:1];
assign y511=x2014[7:1];
assign y767=x3038[7:1];
endmodule